herr talman ! n�got som ocks� beh�vs �r att man i biarritz ser litet l�ngre fram�t .
som de folkvalda vi �r , �r vi �tminstone skyldiga att s�v�l uppmuntra ordf�randeskapet att g�ra framsteg , trots motg�ngarna , som att f�ra vidare de budskap vi f�r fr�n den allm�nna opinionen i v�ra respektive l�nder .
n�r man ser p� h�ndelserna under den senaste tiden tycks mig ocks� fr�gan om bensinpriset s�rskilt anm�rkningsv�rd .
f�r tillf�llet �verv�ger r�det att inkludera en dylik mekanism i artikel 7 .
f�r det andra i �ppenheten f�r medborgarna , som nu vet vilka r�ttigheter de har gentemot dem som till�mpar och skapar europeisk r�tt , och i �ppenheten f�r dem som g�r just detta , skapar eller till�mpar europeisk r�tt .
jag h�ller med honom n�r det g�ller den centrala roll som kommissionen i framtiden skall ha som en garanti f�r det allm�nna gemenskapsintresset .
det �r anledningen till att jag tror att det �r mycket viktigt att ordf�randen i eurogruppen - som vi velat inr�tta - beh�ller hela sin roll i fr�gan .
jag tror f�r min del att det �r just av den anledningen som metoden med konventet �r bra och i h�gsta grad b�r anv�ndas i st�rre utstr�ckning i framtiden .
. ( it ) herr talman , herr r�dsordf�rande , �rade ledam�ter ! jag tackar er f�r den v�nlighet med vilken ni mottog mitt anf�rande och tackar �ven dem som i all v�nskaplighet klandrat mig f�r att jag inte h�llit detta anf�rande tidigare .
vi m�ste arbeta vidare med det f�rst�rkta samarbetet som blivit smidigare och effektivare f�r att uppn� detta resultat : f�rst�rkt samarbete som �r den omedelbara v�gen , den enklaste v�gen f�r att kunna ta steget mot en f�rdjupad integration , vars n�dv�ndighet har bekr�ftats av de m�nga auktoritativa inl�gg som jag har h�rt i dag .
jag f�rklarar h�rmed debatten avslutad .
�ndringsf�rslagen 10 , 11 och 15 �r godtagbara i princip .
denna minskning av parlamentets inflytande �r emellertid godtagbar med tanke p� de ber�rda fr�gornas mycket tekniska natur och kommissionens anstr�ngningar att informera europaparlamentet i god tid om planer p� att utarbeta nya f�rordningar via dess beh�riga st�ndiga kommitt�er .
man vet till exempel att i frankrike varierar siffran f�r skatteinkomster beroende p� om man anv�nder statistik fr�n styrelsen f�r offentliga r�kenskaper eller den fr�n de nationella r�kenskaperna .
en politik i riktning mot en rationell , effektiv och s�ker organisation borde prioritera investeringar i en offentlig europeisk j�rnv�g snarare �n att n�ja sig med att g�ra konkurrensvillkoren mellan v�gtransport�rer enhetliga , vilka framf�r allt �r intresserade av att �ka sina privata vinster .
d� har s�dana bussar visserligen tilltr�de till landet men de kan i praktiken inte n� fram till flera platser .
bet�nkandet st�der r�dets och kommissionens syns�tt och betonar att ett antal reglerande �tg�rder m�ste inf�ras , n�mligen n�r det g�ller pensioner , gr�ns�verskridande prospekt och ett gemenskapspatent .
det sv�raste problemet med denna nya stadga �r inte dess faktiska inneh�ll utan fr�gan om dess juridiska status .
herr talman ! jag r�stade f�r denna stadga , inte minst p� grund av det inflytande som v�r kollega ingo friedrich och professor herzog haft p� inneh�llet i stadgan .
vi menar att stadgan som ett politiskt dokument �r en bra utg�ngspunkt f�r denna helt n�dv�ndiga dialog , som nu skall inledas .
det skulle vara en �verg�ngsl�sning som skulle g�ra det m�jligt att avsluta en stadga med tvingande v�rde .
denna stadga ligger l�ngt hitom den europeiska konventionen om de m�nskliga r�ttigheterna , l�ngt hitom nationella konventioner eller f�rdrag .
. ( fr ) jag r�stade emot ett eventuellt inf�rlivande i f�rdragen av den version av stadgan om de grundl�ggande r�ttigheterna som lagts fram f�r oss .
( a5-0244 / 2000 ) av wiersma om slovakien ( kom ( 1999 ) 511 - c5-0034 / 2000 - 1997 / 2173 ( cos ) ) ;
av den anledningen m�ste det st� klart att det enda som �r v�sentligt �r att fullst�ndigt uppfylla k�penhamnskriterierna .
i det h�nseendet vill jag v�lkomna det arbete som utf�rts av europaparlamentet i form av ett bet�nkande om vart och ett av kandidatl�nderna som inlett f�rhandlingar och ett samlingsbet�nkande fr�n ordf�rande brok , som jag f�r tillf�lle att �terkomma till mer i detalj i mitt inl�gg .
jag t�nker naturligtvis p� den gemensamma jordbrukspolitiken och politiken f�r regional utveckling .
det �r naturligtvis inte uteslutet att kandidatl�nderna tar detta tillf�lle i akt f�r att �nnu en g�ng , - ni talade om det herr talman , - ta upp fr�gan om datum f�r utvidgningen .
utvidgningen �r ett historiskt projekt .
men framg�ngen har inte bara att g�ra med tidpunkten - hur viktig den �n �r .
om de inte f�rverkligas �verallt i europa , d� �ventyras de �verallt .
kapitel p�b�rjas och avslutas i enlighet med den faktiska niv�n p� f�rberedelserna och de faktiska framg�ngarna i f�rhandlingarna .
vad betr�ffar den inre marknaden m�ste vi se till att �verg�ngsfrister b�de tids- och inneh�llsm�ssigt forts�tter att vara s� begr�nsade som m�jligt .
vi beh�ver politiska svar p� politiska fr�gor . de m�ste f�rmedlas p� ett bra s�tt !
t�nk hur vi skulle beh�va l�sa kosovofr�gan , bosnien och hercegovina eller f�rh�llandet till serbien under det kalla krigets dagar .
l�t oss �nd� b�rja debatten med v�r egen befolkning .
vi kommer att kunna och vilja vara med och st�dja allt detta .
mycket av v�r debatt om fruktan inf�r utvidgningen grundar sig p� �verdrifter , men f�r att m�ta de populister som �verdriver , m�ste vi anknyta till en folklig politik genom reflexion .
v�r grupp f�ruts�tter att man i nizza eller omedelbart efter toppm�tet i nizza s�tter ut slutdatum d� medlemsf�rhandlingarna skall slutf�ras .
herr talman ! v�r grupp gruppen europeiska enade v�nstern / nordisk gr�n v�nster h�ller med om m�nga av de tankar och p�st�enden om utvidgningen som ing�r i broks bet�nkande och vi uppskattar den stora insats han har gjort i och med sitt viktiga bet�nkande .
f�r det sj�tte tycker vi att det var ett misstag att i praktiken koppla samman utvidgningen med l�ndernas intr�de i nato .
i likhet med m�nga andra kolleger uppskattade jag i morse mycket det som sades av ordf�rande prodi . jag noterade det som sades av minister moscovici som , med diplomatisk f�rsiktighet , �ven han varnade oss f�r att vi f�r tillf�llet st�r inf�r ett allt annat �n hoppfullt scenario n�r det g�ller de eventuella resultaten under de kommande tv� eller tre m�naderna .
d�rf�r ber jag ministern och kommission�ren att ta h�nsyn till detta n�r det g�ller l�ngden p� inl�ggen .
jag f�r min del drar slutsatsen att vi m�ste tala mer om den , men ocks� tala v�l och b�ttre om den .
jag tror �nd� inte det var en d�lig id� att st�lla fr�gan .
jag vill inte att det d�r skall uppst� n�gra rester , s� som ju varit fallet p� andra omr�den av utlandshj�lpen .
men faktum �r att dagsl�get i dag , den 3 oktober 2000 , �r att jag inte kan s�ga om n�got land i anslutningsprocessen n�r det skall vara moget f�r anslutning .
jag kan ocks� s�ga er varf�r , n�mligen d�rf�r att dessa folk en g�ng f�r alla ville vara p� r�tt sida , dvs. fast f�rankrade i familjen med de demokratiska nationerna .
tack s� mycket f�r ert f�rtydligande , herr kommission�r .
i s� fall har den i mina �gon svikit sitt uppdrag och f�rverkat sitt syfte .
det �r nu som vi kan s�kra gemensamma v�rden och f�rdelar .
f�rest�ll er att en grundl�ggande ekonomisk och samh�llelig omdaningsprocess skulle ha �gt rum i ert eget hemland p� s� kort tid .
hittills har den fortsatt att vara hetluft , herr verheugen , men de faktiska projektansvariga har �nnu inte m�rkt n�got av den .
i dag stabiliserar sig den makroekonomiska situationen .
denna fr�ga kr�ver en s�rskild anstr�ngning och kan , uppskattar jag , inte enbart behandlas som ett biproblem i samband med litauens och polens anslutning .
om vi till exempel betvivlar m�jligheterna f�r medborgarna , f�r arbetstagarna i kandidatl�nderna , att r�ra sig fritt inom europeiska unionen redan fr�n b�rjan , om vi vill f�rv�gra medborgarna i �st denna r�ttighet som utg�r en av unionens grundpelare , s� kommer vi ytterligare att f�rsvaga det folkliga st�det f�r de sv�ra reformer som m�ste genomf�ras inf�r anslutningen .
det gl�der mig att bet�nkandet enh�lligt antogs i utskottet den 14 september .
det handlar f�r min del om - mina kolleger i utskottet f�r utrikesfr�gor , m�nskliga r�ttigheter , gemensam s�kerhet och f�rsvarspolitik har st�tt mig p� denna punkt - att k�penhamnskriterierna , som tjeckerna ocks� har erk�nt - forts�tter att g�lla , och jag �nskar att tjeckerna sj�lva granskar sitt eget r�ttssystem , om s� m�ste vara , sida f�r sida , f�r att unders�ka om det n�gonstans finns n�got som har en diskriminerande karakt�r .
sedan de goda nyheterna , de �verskuggar n�mligen egentligen min kritik .
herr talman , k�ra kolleger ! jag tror att jag kan s�ga att denna rapport , efter att den har debatterats och f�rb�ttrats i utskottet f�r utrikesfr�gor , m�nskliga r�ttigheter , gemensam s�kerhet och f�rsvarspolitik , d�r den fick ett enh�lligt st�d , ganska v�l beskriver och analyserar det nuvarande l�get f�r ungerns anslutning , enligt fr�gans dubbla perspektiv .
det �r en fr�ga som m�ste behandlas seri�st , men i en allm�n ram som omfattar inte bara ungern utan ocks� �vriga kandidatl�nder med denna gamla och os�kra teknik .
misstanken om korruption �r en ytterst destruktiv kraft , som m�ste angripas som ett br�dskande �rende .
i rum�nien har regeringen , med kommission�r verheugens , v�rldsbankens och f�renta nationernas aktiva st�d , gett oss en m�jlighet att uppr�tta goda doktriner och b�sta praxis i regionen .
det handlar om ett kandidatland d�r en tredjedel av territoriet �r ockuperat av den turkiska arm�n sedan 1974 och d�r de grundl�ggande principerna i europeiska unionen p� grund av en ovanligt t�t demarkationslinje inte kan till�mpas p� hela territoriet
europa m�ste bli en ansvarig akt�r n�r det g�ller att l�sa det cypriotiska problemet .
det som �r v�sentligt f�r malta �r det ekonomiska st�det inom ramen f�r anslutningsstrategin och medvetandet om att det st�det f�r malta b�r motsvara de regler som g�ller f�r de andra kandidatl�nderna .
n�r v�l villkoren �r uppfyllda finns det ingen anledning , vare sig f�r kandidatl�nderna eller f�r de nuvarande medlemmarna i eurosamarbetet , att opponera sig mot att kandidatl�nderna g�r in i den tredje etappen av den ekonomiska och monet�ra unionen .
jag �r , om ni s� vill , f�retr�dare f�r en region som f�r tio �r sedan redan utgjorde ett stycke utvidgning �t �ster - ocks� jag levde d� p� andra sidan j�rnrid�n .
i syfte att skapa ett gemensamt informationsomr�de m�ste vi tillsammans f�reta stora anstr�ngningar p� detta omr�de .
�ven tekniskt skiljer sig �st och v�st fortfarande : hos dem finns det fyra internetanslutningar per tusen inv�nare mot sexton hos oss .
i det l�get fick det tidigare �sttyskland massivt st�d med pengar fr�n v�sttyskland , 150 miljarder dm per �r .
under de kommande �ren hotar en avfolkning av landsbygden i �steuropa och �ven ett storskaligt anskaffande av jordbruksmark f�r mekaniserade produktionsintensiva f�retag .
vi bygger upp ett kompendium med direktiv och f�rordningar om fr�gor som har ett tydligt samband med h�lsa , som f�rorening , utsl�pp av radioaktiva och annat farliga �mnen , avfallshantering , vatten- , luft- och markkvalitet , livsmedelss�kerhet samt ansvar f�r nya livsmedel och produkter .
d�rf�r talas det i mitt yttrande inte bara om vad som l�nderna f�r utvidgningen m�ste g�ra , utan �ven om vad europeiska unionen m�ste g�ra .
men nu till de riktiga signalerna .
vi m�ste s�rja f�r att det som nu finns av j�rnv�gsinfrastruktur i central- och �steuropa inte ers�tts med v�gtransporter , s� att man sedan med stor m�da �terigen m�ste f�rs�ka att finna en f�rnuftig l�sning p� det .
detta nej kommer nu att analyseras noga under den n�rmaste tiden .
vi har g�tt igenom texten och har p� ett antal punkter f�rs�kt g�ra vissa saker litet kortare .
man f�r inte offentligt b�rja tvivla p� v�rdet , �ven det omedelbara materiella v�rdet , av den h�r utvidgningen .
om det finns anv�ndning av l�nga �verg�ngssystem p� vissa punkter , l�t oss d� ta i bruk dessa l�nga �verg�ngssystem .
f�r det f�rsta b�r det demokratiska �nskem�let respekteras fr�n ifr�gavarande stater och folk efter anslutningen till eu .
de misstar sig d�rf�r att det �r inte europeiska unionen och dess 80 000 sidor direktiv och f�rordningar som skapar v�lst�nd .
de allt starkare f�rbeh�ll som uttrycks av v�ra befolkningar , liksom danmarks f�rkastande av euron , finns d�r f�r att p�minna oss .
i det yttrande till bet�nkandet brok som jag har varit ansvarig f�r och som budgetutskottet har st�llt sig bakom blir slutsatsen densamma .
perioden h�r inte till de b�sta n�r det g�ller att �gna sig �t utrikespolitik och anklagelserna fr�n de olika partierna kan �ven verka h�gljudda och manipulatoriska .
genom att dela gemenskapens regelverk i tv� delar kunde man � andra sidan s�kerst�lla de nuvarande medlemsl�ndernas integrationsniv� och fr�mja ett intensivare samarbete mellan dem .
jag bes�kte rum�nien i slutet av juli f�r att med egna �gon se hur ett av de st�rsta barnhemmen , som ligger i norra rum�nien , fungerar .
d�rf�r ber vi f�redraganden , kommissionen och r�det att den jordbrukspolitiska delen kompletteras med den fiskeripolitiska delen , exempelvis genom att vi g�r om rubriken " utvidgningens jordbruksaspekter " till " utvidgningens jordbruks- och fiskeriaspekter " .
hellre litet senare och bra �n n�got tidigare och d�ligt .
med cyperns n�ra band till folken i �stra medelhavet , kommer �ns intr�de att st�rka unionens n�rvaro i det viktiga omr�det .
jag st�der f�redragandens �sikt att malta b�r beviljas medlemskap i den f�rsta utvidgningsgruppen och att f�rhandlingarna b�r avslutas f�re utg�ngen av 2001 .
vi �r ocks� ansvariga f�r hur vi f�rmedlar utvidgningen genom ord och handling .
i detta sammanhang handlar det om att skapa opinion f�r utvidgningen .
kommission�r verheugens id� betr�ffande en folkomr�stning om utvidgningen utd�mdes och orsaken �r klar : man kan inte l�ta betalarna besluta om saken .
inf�r den dubbla utmaningen med utvidgningen , som skall g�ra det m�jligt f�r europa att f�rsonas med sig sj�lvt , och den institutionella reformen som skall f�rst�rka demokratin och effektiviteten inom institutionerna , befinner sig europeiska unionen - som s� ofta - vid en viktig v�ndpunkt i sin historia .
jag vill framf�r allt med adress till r�det , som tyv�rr i huvudsak �r fr�nvarande , �nd� uttala n�gra f�rv�ntningar och bet�nkligheter .
en s�dan dialog skulle dessutom bidra till att skapa den administrativa kapacitet som kr�vs f�r en effektiv f�rvaltning av landet , genom att skapa de strukturer som inte finns i dag och minska korruptionen .
malta b�r , liksom de andra mindre medlemsl�nderna , f�retr�das av minst sex ledam�ter .
vi kan inte heller utg� ifr�n att n�got ans�karland naturligt anser sig vara det f�rsta och att utvidgningen inte kan p�b�rjas utan det .
vi hoppas bara att de enorma anstr�ngningar som har gjorts av regeringen den senaste tiden kommer att speglas i kommissionens n�sta rapport .
betr�ffande rum�nien kan man ocks� klarg�ra f�r v�r befolkning att det ligger i v�rt intresse att stabilisera europa .
herr talman ! jag kommer fr�n ett land , sverige , d�r skepticismen mot eu-projektet fortfarande �r ganska stor .
de punkter som utskottet f�r milj� , folkh�lsa och konsumentfr�gor har tillfogat i broks bet�nkande �r steg som �r n�dv�ndiga f�r detta , och en f�ruts�ttning f�r att man skall motverka en stagnation av den europeiska milj�politiken .
sapard-programmet �r en bra m�jlighet till detta , och jag �r mycket positiv till att kommissionen redan har godk�nt sex program .
min grupp har redan meddelat sin �nskan att de f�rsta f�rhandlingarna skall avslutas under �r 2003 , vilket skulle ge en m�jlighet till anslutning i juni 2004 .
den andra minuten vill jag anv�nda till fr�gan om slovenien .
herr talman ! id�n som elmar brok framf�rde h�r i dag betr�ffande ett ees-liknande arrangemang som alternativ f�r de ans�karl�nder som inte uppfyller k�penhamnskriterierna , kommenterades f�rh�llandevis lite .
kandidatl�nderna b�r ocks� uppmuntras att delta i gemenskapens program f�r j�mst�lldhet , i synnerhet ocks� i s�dana som handlar om v�ld mot kvinnor .
men om detta �nd� , trots den cypriotiska regeringens konstruktiva inst�llning , som har erk�nts av alla , visar sig vara om�jligt , p� grund av den turkiska sidans ih�rdiga v�gran , d� anser jag , herr talman , att europeiska unionen inte kan till�ta att cyperns anslutning hindras av den turkiska omedg�rligheten , utan att vi i st�llet omedelbart skall v�lkomna republiken cypern och utn�mna landet till medlem i unionen i avvaktan p� ett framtida , fullst�ndigt deltagande , n�got som f�r �vrigt skedde �ven i fr�ga om en av de grundande medlemsstaterna , vars �rsdag av f�rening vi firar i dag .
justering av protokollet fr�n f�reg�ende sammantr�de
jag anser att det �ven har samband med f�rh�llandet mellan organen att vi ser till att det �ndras !
vi h�ller p� att diskutera en allvarlig fr�ga .
s� �r inte fallet .
detta st�ds i mitt bet�nkande .
mycket av dessa f�rgiftningar eller spridningarna av tunga metaller skedde innan milj�medvetandet var tillr�ckligt och innan man visste vilka effekterna skulle bli .
jag vill l�gga fram ett f�rslag till kommissionen om hur problemet kan hanteras .
de senaste �rens kriser har gjort oss alla mer uppm�rksamma p� detta .
d�rf�r �r vi i europeiska folkpartiets grupp och europademokrater angel�gna om att det skall finnas effektiva kontrollinstrument och vi f�respr�kar , precis som f�redraganden , att kommissionens kontrollexperter oanm�lda i ett n�ra och konstruktivt samarbete med medlemsstaternas kontrollmyndigheter skall kunna utf�ra kontroller p� plats .
vi efterstr�var alla samma sak , och det m�ste ocks� p�pekas h�r .
n�r det g�ller tungmetaller finns det en brist p� konsekvens .
ni m�ste �nd� komma ih�g , mina k�ra kolleger , att eu-institutionernas legitimitet , v�r legitimitet , strikt vilar p� viljan i de nationer som vi har i uppdrag att f�retr�da .
kommissionen har nu f�reslagit att man stryker undantaget f�r foderblandningar och att det finns m�jlighet att fastsl� �tg�rdstr�sklar under de maximalt till�tna gr�nserna vid verklig n�dsituation .
giftrester , f�roreningar , d�lig djurh�llning , d�lig hygien kommer f�rr eller senare att resultera i sjuka djur , och f�ljaktligen ocks� i �kade sjukdomar hos m�nniskorna .
dessa direktiv �r en del av den mest radikala omv�lvningen i gemenskapens hygienbest�mmelser f�r livsmedelss�kerhet sedan minst 25 �r .
jag vill kort ta upp tv� problem vad deklarationen betr�ffar .
jag vill �ven p�peka att det som sker under brottsliga former �r brottsligt !
jordbrukaren m�ste sj�lvklart ers�ttas f�r f�rst�randet av ett f�rorenat och oanv�ndbart spannm�lsparti , liksom man ers�tter till exempel slaktandet av bse-smittade djur .
l�t mig emellertid f�rst ta upp de �ndringsf�rslag som kommissionen inte kan godk�nna .
detta har redan gjorts f�r dioxiner och pcb och man kan f�rv�nta att denna vetenskapliga riskbed�mning finns tillg�nglig som jag sade i oktober .
detta f�rslag �r uppf�ljningen till ett av mina f�rsta �taganden f�r att f�rb�ttra livsmedelss�kerhet och tillhandah�ller ett system f�r att utbyta information p� omr�det djurfoder , med speciell h�nvisning till ett snabbvarningssystem och en r�ttslig grund f�r att kunna inf�ra skydds�tg�rder f�r produkter som framst�llts inom gemenskapen och �ven skyldigheten f�r medlemsstater att ha beredskapsplaner f�r att kunna hantera n�dsituationer som g�ller djurfoder .
i grunddirektivet 95 / 53 fastsl�s redan i artikel 19 att p�f�ljderna f�r icke efterlevnad skall vara proportionerliga och ge en avskr�ckande effekt och n�r det kan bevisas ansvar i civil domstol eller brottsm�lsdomstol g�ller ansvarsskyldighet .
nu har foderblandningsindustrin �ter f�rs�kt att p�verka r�det och stj�lpa den �ppna deklarationen .
vi beh�ver en positivlista med till�tna tillsats- och inneh�lls�mnen f�r djurfoder .
jag anser att insynen i slut�ndan �kar konkurrensen och det uppmuntrar i st�rre utstr�ckning framst�llningen av b�sta t�nkbara blandningar .
d�rf�r anser vi att jordbrukaren skall ha fullst�ndig insyn .
herr talman , herr kommission�r , k�ra kolleger ! efter fr�gan om sammans�ttningen av djurfoder , vilken syftar till att avl�gsna kvicksilver , bly , arsenik , ddt , osv .
vi m�ste skapa realistiska ramvillkor .
herr talman ! f�rslaget som ligger framf�r oss och f�redragandes reaktion p� det �r ett steg i r�tt riktning , men samtidigt kan det inte d�lja den svaga strukturen i kontrollen p� europaniv� .
en omv�nd bevisb�rda , s� som f�resl�s i �ndringsf�rslag 4 , finner jag helt n�dv�ndig med tanke p� de nyss uttalade m�len .
slutligen �r �ndringsf�rslag 6 inte godtagbart d� det inte ligger inom ramen f�r detta direktiv .
det �r n�r vi skall r�sta om dessa punkter som jag kommer att fr�ga om det finns n�gra inv�ndningar mot att de f�rs in efter punkt 1 .
( kammaren godk�nde att det muntliga �ndringsf�rslaget tas upp till omr�stning . ) ( parlamentet antog resolutionen .
( parlamentet antog resolutionen . )
f�r det andra att kandidatl�nderna forts�tter med sin positiva utveckling f�r att uppfylla k�penhamnskriterierna och mot ett fullst�ndigt genomf�rande av gemenskapens regelverk f�re anslutningen .
punkt 65 vittnar ocks� om bryssels hegemoniska och likriktande vilja , eftersom det f�rklaras att icke-diskrimineringsklausulen i artikel 13 i eg-f�rdraget �r en del av gemenskapens regelverk och man h�vdar att " lagstiftning som grundar sig p� denna till fullo b�r inf�rlivas i l�nderna i central- och �steuropa " .
f�r att �terkomma till de finansiella aspekterna : det verkar vara n�dv�ndigt att studera de finansiella �terverkningarna av att det tillkommer ett s� stort antal nya medlemsstater , innan den nuvarande budgetperioden har l�pt ut �r 2006 .
n�r kandidatl�nderna ansluter sig till eu skall de behandlas likv�rdigt med alla andra medlemsl�nder inom eu . vi kan under inga omst�ndigheter acceptera att nya medlemsstater behandlas som andra klassens medlemmar .
det motsatta f�rh�llandet skulle orsaka splittring inom jordbruket och utg�ra en fara f�r den sociala utvecklingen i hela europas lantliga struktur .
i detta bet�nkande f�resl�s i realiteten en utvidgning av en ekonomisk marknad .
riskerna �r att unionen urvattnas politiskt och att social dumping blir vanligt , och slutligen att det europeiska projektet begr�nsas till en stor marknad och ett omr�de med fri konkurrens .
p� pappret har mycket uppn�tts in puncto likabehandling och lika m�jligheter f�r kvinnor och m�n . men hur ser det ut i praktiken ?
. ( fr ) europeiska unionens utvidgning till tio l�nder i �steuropa samt malta och cypern �r ett stort projekt .
f�r det andra : utvidgningen medf�r oundvikligen att europeiska unionen m�ste se �ver sina ekonomiska planer som uppr�ttades och fastst�lldes innan utvidgningen var p�t�nkt .
herr talman ! det �r mig ett stort n�je att meddela att jag r�stade f�r �tg�rden om estlands ans�kan om medlemskap i europeiska unionen .
jag konstaterar att lettland g�r framsteg f�r att uppfylla b�de k�penhamnskriterierna och f�r att uppfylla skyldigheterna i fr�ga om gemenskapens regelverk .
jag konstaterar att litauen g�r goda framsteg att uppfylla b�de k�penhamnskriterierna och skyldigheterna som g�ller gemenskapens regelverk .
polen respekterar dessutom fullt ut de m�nskliga r�ttigheterna och de grundl�ggande friheterna .
polen har alltf�r l�nge betraktats som sina hotfulla grannars fr�msta slagf�lt , f�r vilka en annektering av polen alltid har varit den f�rsta punkten p� deras expansionistiska program ; det har betraktats som en ofrivillig scen f�r historiens mest avskyv�rda tragedier och sedan , under flera decennier , som ett land vilket �verl�ts till f�rtrycket under en totalit�r regim , som med uppmuntran av v�r medbrottsliga tystnad trodde sig ha f�tt bukt med landets legendariska motst�ndsanda . men polen har aldrig upph�rt att med stor kraft illustrera v�rden som frihet , mod och oberoende - allt det som utg�r grunden f�r de gemensamma v�rderingar p� vilka v�rt politiska europabygge f�rv�ntas vila .
om tjeckien forts�tter sitt framg�ngsrika arbete och europeiska unionen anpassar sin institutionella struktur och politik f�r att klara utvidgningen ser jag inget hinder f�r tjeckien att kunna ansluta sig till unionen .
" till republiken ungern allts� .
om bulgarien forts�tter att utvecklas positivt och europeiska unionen anpassar sin institutionella struktur och politik f�r att klara utvidgningen ser jag inget hinder f�r bulgarien att kunna ansluta sig till unionen .
jag hoppas att slovenien kommer att finnas i den f�rsta gruppen av nya medlemsl�nder .
fr�gan om flyktingarnas �terv�ndande och om bos�ttningarna p� cypern tas upp .
det �r f�r �vrigt kontentan av slutsatserna fr�n europeiska r�dets m�te i helsingfors , d�r man �ntligen bekr�ftade att en l�sning p� cypernfr�gan inte utg�r ett " n�dv�ndigt villkor " f�r ett eu-medlemskap .
vi hoppas att utsikten om ett tidigt medlemskap i eu och underl�ttandet av kontakter med hj�lp av samlevnadsprojekt fr�n gr�srotsniv� och upp�t som eu lovat att st�tta och finansiera kan ge en positiv input till l�sningen av " cypernfr�gan " .
det f�rekommer avsiktliga brott mot sanit�ra f�reskrifter , straffr�ttsliga best�mmelser och t.o.m. moraliska regler , eftersom naturens lagar f�rfalskas och arter och djurens fysiologi inte respekteras , utan att det g�rs n�gra som helst kontroller , utformas l�mpliga regler och utf�rdas motiverade straff .
vi m�ste faktiskt visa vaksamhet p� det h�r omr�det , eftersom djurfoder utg�r den f�rsta l�nken i livsmedelskedjan .
mot bakgrund av det f�rflutna och dagens ekonomiska f�rbindelser mellan de utvecklade stormakterna och asiens fattiga l�nder , �r det i b�sta fall en from �nskan att tala om " j�mb�rdiga partner " f�r framtiden , men mera troligt �r det ett s�tt att med pseudo-demokratiska och pseudo-humanit�ra fraser d�lja det faktum att f�rbindelserna grundas p� exploatering .
jag vill p�peka f�r ledam�terna att r�dets arbetsgrupp var enh�lligt �verens om att rekommendera r�det att kommitt�n i handlingsprogrammet b�r �ndras till blandad kommitt� , en kombination av f�rvaltnings- och r�dgivande f�rfaranden och d�rigenom �ka de enskilda medlemsstaternas befogenheter .
jag f�rst�r deras oro men jag har f�rs�kringar fr�n kommissionen att frist�ende organisationer fortfarande kommer att kunna ans�ka om bidrag f�r detta och andra program och initiativ som kommissionen organiserar .
d�rf�r �r det absolut n�dv�ndigt att de grupper som omn�mns i artikel 13 skyddas effektivt fr�n diskriminering .
f�r det fj�rde : arbetsmarknadens parters deltagande .
det har fullt klargjorts f�r mig hur mycket vi beh�ver ett s�dant mot bakgrund av utfr�gningarna om artikel 13 .
principiell av det sk�let att likabehandling �r en grundl�ggande r�ttighet , vilken som s�dan �r en av de grunder som europeiska unionen vilar p� .
den budgetsp�nning som finns i utgiftsomr�de 3 , d�r detta och andra program h�r hemma , �r ingen hemlighet f�r n�gon , k�ra kolleger .
undantag med en annorlunda behandling som kan etableras av ideologiska och religi�sa sk�l , eller av �lderssk�l , m�ste f�rena den r�tt vissa offentliga eller privata organisationer �tnjuter med en noggrann respekt f�r lika behandling .
betr�ffande de n�rmare detaljerna i bet�nkandet vill jag tacka herr mann som godtog de flesta synpunkterna fr�n utskottet f�r industrifr�gor , i synnerhet dem som g�llde m�ngsidig diskriminering - som i fallet kvinnor , som uts�tts f�r annan diskriminering .
vi h�rde dem f�r flera �r sedan betr�ffande lika l�n f�r kvinnor , vi h�rde dem n�r vi lagstiftade om j�mlikhet , f�rb�ttrad mammaledighet , vi h�rde dem i samband med rasdirektivet f�re sommaren s� vi m�ste obekymrat g� vidare .
den ber�r fr�gan om m�ngfald . det �r m�nga som inser hur viktigt detta �r f�r att v�r demokrati skall fungera v�l .
jag skulle f�r �vrigt ocks� vilja ta tillf�llet i akt f�r att �ven gratulera kollega cashman , f�r direktiv �r viktiga , men handlingsprogram f�r att st�dja dem �r naturligtvis ocks� oumb�rliga .
herr talman , fru kommission�r , k�ra kolleger ! b�da f�redraganden har �stadkommit ett fantastiskt arbete som jag vill tacka f�r som f�retr�dare f�r min grupp .
d�rf�r �r vi mycket tveksamma till denna punkt och ber att kommissionen , n�r den skall kontrollera hur dessa medel anv�nds , ser upp s� att inte turkiet l�tsas utrota eller bek�mpa diskrimineringen av br�drafolket utan att egentligen alls avskaffa den grundl�ggande diskrimineringen som verkligen �r den som ligger till grund f�r m�nga olyckor f�r v�rt europa .
personalen , s�v�l i chefsst�llning som underordnade , skapar gemensamt formen f�r detta .
jag tror att vi d�rigenom bara skapar st�rre os�kerhet , eftersom vi inte l�ngre vet , vem som kan st�djas i enlighet med kommissionens program .
herr talman , fru kommission�r ! v�r grupp har bed�mt b�da bet�nkandena positivt och vill s�rskilt understryka hur koncentrerade alla �r p� behovet att utvidga programmets till�mpningsomr�de genom en rad �ndringsf�rslag - som faktiskt har visat p� m�nga nya former av diskriminering - f�r att f�rs�ka s�kerst�lla att alla m�nniskor behandlas likv�rdigt oberoende av k�n , ras , etniskt ursprung , religion , personlig �vertygelse , �lder och sexuell l�ggning .
syftet med detta arbete grundat p� artikel 13 �r att g�ra j�mlikhet till en realitet genom att ta bort det leende ansikte som s� ofta d�ljer f�rdomar och tr�ngsynthet , framf�r allt p� arbetsplatsen .
artikel 5 , i dess nuvarande form , har kritiserats f�r att den verkar f�rsvara det som den syftar till att bek�mpa .
men sedan 40 �r tillbaka finns det ocks� texter som tv�rtom vilar p� diskriminering .
generellt sett �r jag positiv till att man betonar vikten av att utveckla och ut�ka de kulturella aspekterna n�r det g�ller diskriminering , jag tror rent av att diskrimineringen kan �vervinnas genom en kultur av icke-diskriminering , genom att ge aktuell och l�ttillg�nglig information till alla medborgare i alla medlemsstaterna .
herr talman , fru kommission�r , �rade ledam�ter ! som bekant finns det fortfarande mycket diskriminering i europeiska unionen , fr�mst n�r det g�ller syssels�ttning och yrkesverksamhet , trots f�rbuden enligt artikel 13 i f�rdraget om europeiska unionen .
jag v�lkomnar detta direktiv som det allra f�rsta eu-lag som i hela europa inf�r r�ttigheter f�r v�ra 37 miljoner medborgare med funktionshinder ett slut p� att via bakd�rren lagstifta om handikappades r�ttigheter och en hyllning till handikappr�relsen som har drivit kampanjer f�r att uppn� denna dag .
detta �r vad som skiljer vissa b�nkar fr�n andra .
insatsen kommer annars inte att bli en framg�ng i verkliga livet .
slutligen m�ste europaparlamentet h�llas informerat och kammarens bet�nkanden och yttranden skall beaktas . vi b�r ocks� framh�va vikten av att icke-statliga organisationer och f�reningar verkligen kommer med sina �sikter och deltar - och de b�r f� n�dv�ndiga medel - f�r de �r helt klart nyckelakt�rer f�r att de antagna �tg�rderna skall n� framg�ng .
den best�mmelse som s�ger att det kan g�ras undantag till begreppet yrkesmeriter - ett mycket viktigt och avg�rande begrepp - med h�nvisning till en religion , den �r inte godtagbar f�r mig .
v�r gemensamma civilisation bekr�ftar sin storhet genom respekten f�r det �ppna , toleranta och liberala samh�llet och genom dess m�ngkulturella politik som inkluderar alla .
. ( en ) som ni k�nner till f�reslog kommissionen i november ett stort paket baserat p� artikel 13 med tv� direktiv och ett program .
kort sagt jag kan d�rf�r varken som f�rslag eller i andan godk�nna �ndringsf�rslagen 1 , 2 , 7 , 8 , 10 , 11 , 13 , 18 , 21 , 41-45 , 47 , 50 , 58 , 59 , 62 , 64 , 65 , 66 och 67 .
med dessa tv� till�gg anser jag att f�rslagets r�ckvidd blir tydlig .
jag vill g�rna i detalj ta upp de �ndringsf�rslag som jag inte kan godk�nna eftersom de skapar politiska och r�ttsliga sv�righeter .
detta direktiv m�ste vara en del av det sociala regelverket i ans�karl�nderna .
dessutom k�ar icke eu-l�nder f�r att ansluta sig till koden .
jag gl�der mig av hela mitt hj�rta �ver denna utveckling .
jag uppmanar alla andra regeringar att g�ra detsamma .
d�rf�r mots�tter vi oss ocks� de �ndringsf�rslag som ingivits av v�ra kolleger , vilka kr�ver en allm�n nedrustning p� internationell niv� och att europeiska unionen b�r vara den som visar v�gen .
spridningen av l�tta vapen forts�tter att vara orov�ckande , �ven i v�rt n�romr�de , till exempel p� balkan .
sverige anser inte att verksamheten inom gusp kan beskrivas som f�rsvarspolitik , eftersom den inte inneb�r n�gon gemensam f�rsvarsf�rpliktelse motsvarande natos paragraf 5 .
i eu : s uppf�randekod fastsl�s en upps�ttning av utf�rliga principer f�r konventionell vapenexport .
europeiska unionen har f�rbundit sig att bek�mpa den destabiliserande effekten av f�r stora m�ngder handeldvapen i m�nga delar av v�rlden .
jag vill �terigen tacka f�redraganden f�r hans utm�rkta bet�nkande , som inneh�ller en stor m�ngd anv�ndbara anvisningar om hur vi skall utvecklas v�r politik p� detta ytterst viktiga omr�de .
dit kan vi n� genom att till�mpa de kriterier som anv�nds f�r att fastst�lla detta merv�rde , med sikte p� rangordning och uteslutning .
men hittills har det inte n�dv�ndigtvis f�rekommit en rangordning , och inte heller faktorer f�r uteslutning .
herr talman ! jag skulle vilja tacka kommission�ren f�r hans inledning , men jag har �nd� ett par fr�gor .
ni som har erfarenhet kanske s�ger att det redan har p�pekats flera g�nger .
f�r att till sist svara pi�trasanta vill jag tacka honom f�r hans anf�rande och konstruktiva vilja .
herr kommission�r ! jag tackar er f�r er n�rvaro h�r och f�r det meddelande som ni har redogjort f�r .
den socioekonomiska forskningen har helt klart sin plats .
jag vill ocks� s�ga att jag �r bekymrad �ver den mycket l�ga niv� p� sammanh�llningsfondens �tagandebemyndiganden som g�llde i slutet av augusti - endast 16 procent , fru ledamot - samt bekr�fta , �ven om utvecklingen har g�tt i r�tt riktning sedan slutet av augusti , mina farh�gor som jag den 11 september delgav utskottet f�r regionalpolitik , transport och turism .
men jag tror , herr kommission�r , urs�kta att jag s�ger det , att ni inte �r s� v�linformerad .
kan ni ge oss siffrorna f�r spanien och grekland ?
det f�rslaget st�tte dock p� massivt motst�nd fr�n vissa medlemsstater .
om br�nslekostnaderna i ett f�retag som detta �r mer �n dubbla mot dem f�r multinationella f�retag med andra baser p� andra h�ll i skottland som kan l�gga in anbud f�r samma kontrakt , snedvrider detta uppenbarligen konkurrensen till nackdel f�r avsides bel�gna samh�llen .
mot bakgrund av gemenskapens �tagande f�r att uppfylla �tagandena fr�n kyoto undrar jag om kommission�ren skulle godk�nna att det b�sta s�ttet att g�ra detta �r genom h�gre br�nsleskatter i motsats till att h�ja andra transportkostnader .
om kommissionen inte har instrument f�r att p�verka niv�erna p� punktskatter i medlemsstaterna och om det enligt konkurrensreglerna inte �r till�tet att gynna vissa industrier d� skulle det v�l , n�r en region blir lidande p� grund av att den ligger i ett yttre eller avl�gset omr�de , vara fr�ga om utj�mnande insatser inte om att ge n�gra speciella f�rdelar om det fanns n�gra skillnader i de till�tna punktskatterna under dessa speciella och s�rskilda omst�ndigheter ?
det finns emellertid inga specifikt reserverade belopp f�r minoritetsspr�k inom ramen f�r dessa aktiviteter , vilket inte hindrar att dessa program anv�nds f�r dessa syften .
. ( en ) jag skall besvara fr�gorna fr�n herr sacr�deus och fru theorin om samma �mne samtidigt .
jag undrar om �rendet har bollats fram och tillbaka mellan olika eu-kommission�rer utan att n�gon i slut�ndan tagit ett verkligt ansvar f�r fr�gan .
varje �r tvingas �ver 1 miljon barn in i barnprostitution .
betr�ffande kompensation anser medlemsstaterna och kommissionen att offentliga myndigheter och privata , ekonomiska akt�rer sj�lva skall b�ra kostnaderna f�r omst�llningen inom sina respektive omr�den .
. ( en ) herr talman ! helt kort , elva l�nder har godk�nt euron .
j�garf�rbunden skall spela en viktig roll f�r att s�kerst�lla att j�gare har kompetens att g�ra en s�dan bed�mning .
vad g�ller frankrike v�ntar kommissionen p� information om vilka �tg�rder som vidtagits av de ber�rda myndigheterna r�rande n�gra av rekommendationerna i fvo-rapporten , bland annat om vilken �tg�rd som vidtagits f�r att se till att f�rdplaner anv�nds och undertecknas ordentligt .
jag skulle vilja att kommission�ren ber�ttade lite mer om den speciella fr�gan om �vertr�delsef�rfaranden mot italien .
kommissionens enheter utarbetar just nu ett f�rslag till kommissionens direktiv som r�r dessa fr�gor , d�ribland bomullsfr�n .
. ( en ) detta �r en fr�ga som i sj�lva verket faller inom min kollegas , herr liikanen , ansvarsomr�de .
herr talman ! jag tackar kommission�ren f�r den informationen och f�r n�gra bevis p� framsteg i granskningen av denna fr�ga .
den spanska regeringschefen - aznar - kommer i oktober att g�ra ett officiellt bes�k i iran .
jag f�renar mig med den �rade ledamoten och uttrycker min beundran f�r aung san suu kyi och hennes partikamrater i nld .
levnadsf�rh�llandena f�r folket i burma , p� grund av den hemska regering som drabbat dem , �r sv�ra nog som de �r , och jag skulle inte vilja g�ra n�got som f�rv�rrade dessa levnadsf�rh�llanden .
jag hoppas att vi skall kunna forts�tta att ge humanit�r hj�lp till dem , men det som uppenbarligen �r mest viktigt - det skulle uppmuntra dem att �terv�nda fr�n bangladesh och fr�n andra l�nder i regionen - det som �r mest viktigt �r att det blir en politisk �verenskommelse d�r dessa r�ttigheter erk�nns liksom r�ttigheterna f�r dem som blev demokratiskt valda f�r �ver tio �r sedan men som generalerna drev undan .
n�r jag bes�kte kosovo h�romdagen gjorde det starkt intryck p� mig att m�nniskor talade om f�r mig att den f�rsta etappen av valkampanjen hade genomf�rts ytterst professionellt .
jag f�rklarar h�rmed fr�gestunden avslutad .
det b�r ske grundliga multilaterala samr�d innan ett land beviljar en licens som ett annat land har avslagit .
den teknik och expertis som finns tillg�nglig b�r anv�ndas till n�got konstruktivt i samh�llet , n�got som skall gagna m�nniskor snarare �n n�got som skall f�rinta och f�rst�ra m�nniskor .
kontrollmekanismen m�ste framf�r allt utstr�ckas f�r att omfatta l�tta vapen och finkalibriga vapen som anv�nds i m�nga regionala och etniska konflikter i v�rlden , och som ofta riktas mot civil och milit�r personal fr�n eu-l�nderna .
herr talman ! jag �r glad att s� m�nga personer fr�n allm�nheten h�r i dag f�r alla d�r uppe kan se finns det mycket f� personer n�rvarande h�r nere vid denna tid p� kv�llen .
medan utskottet �r positivt till det v�sentliga i kommissionens f�rslag finns i mitt bet�nkande ett antal �ndringar som m�ste g�ras f�r att f� f�rslaget om �tskilda befogenheter att fungera .
ett av de problem som parlamentet har haft under senare �r �r bristen p� standardiserad information om budgetkontroll fr�n institutionerna .
" utmaningen f�r kommissionen kommer att vara att �vertyga parlamentet att den kan skapa denna s�kerhet .
resultat : den nya mannen i ledningen kommer visserligen utifr�n , men han fastnar genast i f�llan av en redan f�rdiginstallerad apparat .
det finns enligt v�r uppfattning en dissonans i bet�nkandet , men min grupp �r inte enig om detta , och det g�ller fr�gan om internkontrollen enbart skall inr�ttas f�r kommissionen , r�det och parlamentet eller �ven f�r de mindre institutionerna ?
det f�rv�ntar vi oss mycket av .
herr talman ! jag vill inleda mitt inl�gg med att gratulera hulten till detta s� v�l genomf�rda bet�nkande som fick ett enh�lligt st�d av kollegerna i budgetkontrollutskottet .
enbart det faktum att det kan verka som att det inte l�ngre f�religger ett oberoende , borde f� oss att �ter betrakta den funktionen separat .
jag vill d�rf�r �ter po�ngtera att vi har utvecklat ett mycket exakt f�rfarande f�r att unders�ka om de enskilda generaldirektoraten som i forts�ttningen kommer att vara ansvariga f�r dessa f�rhandskontroller �r i st�nd till detta .
jag vill bland annat p�minna om att det i artikel 22.2 i direktivet , uttryckligen st�r att alla medlemsstater skall vidta l�mpliga �tg�rder f�r att tv-bolagens uts�ndningar inte skall inneh�lla n�gra program som kan skada minder�rigas fysiska , mentala eller moraliska utveckling , s�rskilt program som inneh�ller pornografiska scener eller on�digt v�ld .
vi vill inte byta ut den som g�r n�got gott i nationerna , men vill p� gemenskapsniv� inf�ra gemensamma kriterier och minimikrav , f�resl� best�mmelser som hj�lper m�nniskor i de olika l�nderna att verkligen oms�tta uppgiften att skydda de minder�riga i praktiken .
de problemen g�r inte att komma �t med hj�lp av tekniska anordningar f�r kontroll av tv-s�ndningar .
kommissionens ordf�rande , romano prodi , n�mnde i sitt stora , fina tal i g�r , att det med h�nsyn till eu : s politiska legitimitet i framtiden kommer att bli n�dv�ndigt att utarbeta en katalog �ver vilka fr�gor som eu skall syssla med , och vilka fr�gor medlemsstaterna skall syssla med .
herr talman , fru kommission�r ! nyttjandet av och tillg�ngen till tv , tryckt material och nya medier h�r till v�ra barns vardag och �r f�r dem en sj�lvklarhet .
herr talman , fru kommission�r , k�ra kolleger ! det var en s�ndag kv�ll f�r tv� veckor sedan i s�dra frankrike , n�r johan 17 �r och robert 16 �r d�dade romain , deras barndomskompis , med ett eldvapen och ett basebolltr� , utan anledning , utan syfte - som p� tv .
barnen kommer att kunna hantera dessa filtersystem b�ttre �n vi , och det mycket snabbt .
kommissionen skall beakta denna uppmaning , eftersom ni vet att vi �r 2002 skall l�gga fram direktivet " television utan gr�nser " p� nytt , f�r att g�ra en �versyn .
vi m�ste se till att erfarenheten hos ungdomar - studenter och �vriga som finns i utbildningsv�rlden - �r positiva .
jag hoppas d�rf�r att vi �ntligen skall finna en definitiv l�sning s� att r�rligheten i europeiska unionen - f�r studerande , m�nniskor som yrkesutbildar sig , unga frivilligarbetare , l�rare och yrkesl�rare - blir en fj�der i hatten f�r europeiska unionen och s� att vi kan undvika den paradox som s�ger att det �r l�ttare f�r varor , kapital och tj�nster att r�ra sig i europeiska unionen �n f�r de europeiska medborgarna sj�lva .
herr talman ! jag beklagar att ungdomar h�rigenom hindras att skaffa sig erfarenhet , studieerfarenhet , arbetserfarenhet eller annan erfarenhet , i en annan medlemsstat .
jag hoppas att de viktiga �ndringsf�rslag som godk�nts av utskottet f�r kultur , ungdomsfr�gor , utbildning , medier och idrott f�r det positiva gensvar av r�det som de f�rtj�nar och att lagstiftningen snabbt kan tr�da i kraft .
fri r�rlighet f�r personer , varor , tj�nster och kapital finns bekr�ftad i v�ra f�rdrag och �nd� v�gras unga m�nniskor , som �r europeiska unionens framtid och kanske har mindre f�rdomar �n n�gra av oss vuxna , m�jligheter p� grund av byr�kratiska hinder som finns i deras v�g .
men det universitet som inte erk�nner utbildningar b�r f� sina bidrag indragna .
just d�rf�r �r jag fortfarande f�rv�nad �ver att det f�religger s� m�nga hinder f�r en �kad r�rlighet och flexibilitet i europa .
s� trots de problem som kvarst�r , och jag k�nner till dem , �r dessa program positiva och medf�r n�got till befolkningen .
tack s� mycket , kommission�r reding .
den 6 juli i leipzig framf�rde ni en v�djan om en fram�tblickande vision av europa , grundad p� ett f�rfattningsprojekt .
n�r det g�ller att uppn� dem , i sin helhet och i tid , pr�vas v�r f�rm�ga att konsekvent genomf�ra det vi s�ger oss vilja g�ra .
och �nd� ligger europa vid medelhavet !
jag kommer i dag att tala om ett j�mlikt deltagande av kvinnor och m�n p� samtliga samh�llsomr�den .
�tg�rdsprogrammet fr�n peking och de senaste rekommendationerna i juni fr�n det s�rskilda sammantr�det i fn : s generalf�rsamling om peking + 5 g�r i samma riktning .
jag vill ge tv� exempel : r�det f�r utbildning vad g�ller fr�gan om manliga och kvinnliga studerandes r�rlighet samt manliga och kvinnliga l�rares r�rlighet , eftersom vi har blivit medvetna om att det finns stora olikheter i fr�ga om r�rlighet , samt r�det f�r den inre marknaden , konsumentfr�gor och turism vad g�ller fr�gan om utveckling av elektronisk handel f�r att g�ra den tillg�nglig f�r alla m�n och kvinnor , eftersom vi vet att ocks� h�r finns det olikheter mellan m�n och kvinnor vad g�ller elektronisk handel .
den f�rsta artikeln �gnas �t den allm�nna principen f�r j�mst�lldhet inf�r lagen f�r alla m�nniskor .
jag vill d�rf�r g�rna v�dja till r�dets ordf�rande , b�de den nuvarande och den kommande , och kommission�ren om att vara uppm�rksamma p� denna aspekt , d�rf�r jag tror att det �r helt grundl�ggande f�r v�rt arbete att vi g�r en mycket stor insats p� detta omr�de .
om vi nu tar en titt p� j�mlikhetspolitiken s� tycker jag det verkar , nu n�r vi sitter h�r allihop och det �r huvudsakligen kvinnor som sitter h�r och som deltar i diskussionen , som om vi alla naturligtvis g�r v�rt allra b�sta , men att vi ocks� �r medvetna om att den europeiska j�mlikhetspolitiken riskerar att f�rlora sin slagkraft .
n�gra problemomr�den : kvinnor �r ofta dubbelarbetande , arbetsl�sheten �r h�gre bland kvinnor , barnomsorgen har f�rs�mrats , det finns f�r f� kvinnor i beslutande st�llning , kvinnov�ldet �kar i m�nga kandidatl�nder , och fler kandidatl�nder �r centrum f�r den �kande kvinnohandeln .
pery talade om vikten av att f�rena arbete och familjeliv .
vi m�ste se till att det som beslutas i strasbourg �r ett verkligt framsteg .
i st�llet f�r att v�nda sig till alla , delar vi upp i fack , efter minoritet och efter folkgrupp .
andra ledam�ter av parlamentet var tvungna att ta till pennan f�r att tillr�ttal�gga . polen tackade dem f�r det f�r �vrigt .
barnuppfostran , s�rskilt �verf�ringen av normer och v�rden �r livsviktigt f�r v�rt samh�lle .
f�r det f�rsta f�r att f�rb�ttra de befintliga direktiven , till exempel om likabehandling av m�n och kvinnor i f�retags- eller yrkesbaserade system f�r social trygghet .
jag var f�redragande i peking och vice f�redragande i new york .
jag st�der beg�ran i detta bet�nkande fr�n utskottet f�r kvinnors r�ttigheter och j�mst�lldhetsfr�gor om en omfattande kvinnounders�kning i eu och ans�karl�nderna som en inledning till ett framtida arbete .
dagligen konstaterar vi , �ven efter folkomr�stningen i danmark nyligen , att detta �r ett omr�de d�r vi m�ste g�ra n�got . vi anser det ocks� n�dv�ndigt att kvinnorna , b�de kvalitativt och kvantitativt , �r politiskt aktiva i de olika medlemsstaterna och , om m�jligt , i europas olika regioner , s� att de medverkar i kommissionens initiativ och program , f�r jag anser att det r�der stor brist p� information mellan kvinnor i allm�nhet och de organiserade kvinnogrupperna , men ocks� en obalans i fr�ga om aktivt politiskt deltagande mellan olika omr�den i europa .
detta �r allts� en oerh�rt viktig fr�ga f�r oss att ta tag i .
herr talman ! jag vill uttrycka min uppskattning �ver perys n�rvaro h�r i kammaren liksom �ver kommission�r diamantopoulous n�rvaro .
. ( fr ) herr talman , jag kommer inte att svara var och en enskilt , utom torres marques , eftersom hennes fr�ga verkligen �r alltf�r direkt och personlig .
den fj�rde fr�gan : framtidsfr�gorna .
f�r det andra , d�rf�r att de ger en m�jlighet till j�mf�relser mellan medlemsstaterna , men ocks� en j�mf�rande utv�rdering av utvecklingen inom europeiska unionen som helhet .
jag skulle �nnu en g�ng vilja tacka dybkjaer f�r jag anser att hon lagt ner ett utomordentligt stort arbete p� sitt bet�nkande , som kommer att vara till stor nytta f�r oss i v�r n�sta rapport , och jag vill speciellt tacka det franska ordf�randeskapet och pery f�r att de under denna tid gripit sig an j�mst�lldhetsfr�gorna med s� stor energi .
tre av dessa - �ndringsf�rslag 4 , 5 och 7 - g�llde kommitt�f�rfarandet .
utskottet f�r r�ttsliga fr�gor och den inre marknaden har - som f�redragande p�pekade - godtagit det resonemanget och d�rf�r avst�tt fr�n att l�gga fram �ndringsf�rslagen p� nytt .
om vi d�rf�r medger , som r�det och kommissionen sade , att det �ndringsf�rslaget inte �r l�mpligt i det h�r fallet , vill jag �ter passa p� att p�minna om att f�rfarandena f�r kontroll av import till europeiska unionen inte fungerar , att bedr�gerier sker , och att dessa bedr�gerier inte bara �r negativa f�r gemenskapens skattebetalare utan ocks� f�r den inre marknadens funktion och dessutom f�r lojaliteten gentemot tredje land .
det �ppnar v�gen f�r en viktig reform av de ekonomiska tullsystemen , om vilka parlamentet f�rresten skall f� detaljerad information om f�r godk�nnande under de kommande m�naderna .
i g�r f�r�ndrades hela st�ndpunkten i och med den st�ndpunkt kommissionen redovisade i samband med den r�ttsliga grunden .
herr ordf�rande ! det �r en stor gl�dje f�r oss att v�lkomna er till europaparlamentet och vi hoppas att ni kommer att trivas under ert bes�k .
( parlamentet antog resolutionen . )
de europeiska medborgerliga r�ttigheterna verkar inte v�ga s�rskilt tungt i situationen .
ut�ver en symbol �r det en motivation och en motor f�r tillh�righet i den kultur och den modell f�r europeiskt samh�lle som vi g�r anspr�k p� .
herr talman ! jag r�stade f�r cashmanbet�nkandet , f�r ordf�randen f�r pension�rsf�reningen i den kommun d�r jag bor - curno i provinsen bergamo i italien - sade till mig : " vi har inga som helst m�jligheter att f�rsvara de �ldres intressen .
oavsett sina olika st�ndpunkter i �vrigt har de visat att , n�r ett �ndringsf�rslag �r riktigt , s� st�der de det , oavsett vem l�gger fram det .
den best�mmelse enligt vilken begreppet om v�sentliga och avg�rande yrkesm�ssiga krav kan ligga till grund f�r religionsgrundade undantag riskerar att bli f�rem�l f�r en bred tolkning .
parallellt m�jligg�r det �ndringsf�rslag genom vilket undantaget fr�n principen om icke-diskriminering breddas till att omfatta religi�sa organisationers sociala verksamheter i vid mening , om det g�ller diskriminering som enbart grundas p� religi�sa �vertygelser och inte n�got annat sk�l , s� att dessa strukturers specifika pr�gel och annorlunda insats st�rks i f�rh�llande till offentliga eller privata tj�nster .
vissa , s�kert v�lmenta , �ndringsf�rslag som vi fick ta del av f�r en att undra om m�nniskan alltid l�ter f�rnuftet segra .
. ( en ) eplp ( european parliamentary labour party ) har r�stat f�r mann-bet�nkandet om likabehandling i arbetslivet , eftersom eplp p� ett best�mt s�tt tar fasta p� principen om bek�mpning av or�ttvis diskriminering och att vi kan uppvisa ett brett st�d f�r de �vergripande m�len bakom detta f�rslag .
vi hyser bet�nkligheter n�r det r�r inbegripandet av h�lso- och sjukv�rd , social trygghet och bist�nd , eftersom det finns avsev�rda nationella skillnader n�r det g�ller hur dessa fr�gor hanteras , och om de utg�r en del av f�rh�llandet mellan arbetstagaren och arbetsgivaren .
" tack vare agerandet av en " ringare " och het de vises kommitt� har korruptionen kunnat f�rd�mas .
vi i europa , tillsammans med v�ra kolleger �ver hela v�rlden , m�ste se till att g�ngna tiders misstag och girighet inte upprepas .
bet�nkandet ser vapenexportkontroll huvudsakligen som en metod att undvika obekv�ma situationer f�r europas milit�rindustri och inte som en s�tt att �stadkomma nedrustning och fred .
. det �r bra att europeiska unionen vill genomf�ra en uppf�randekod f�r en restriktiv vapenexport .
bet�nkande ( a5-0258 / 2000 ) av angelilli
jag vill p�minna er om att med st�d av best�mmelserna i artikel 22c.2 i direktivet om television utan gr�nser ( direktiv 97 / 36 / eg av den 30 juni 1997 om �ndring av direktiv 89 / 552 / eg ) var kommissionen skyldig att g�ra en unders�kning om eventuella f�r- och nackdelar med �tg�rder i syfte att l�tta p� f�r�ldrarnas eller l�rarnas kontroll av de program som minder�riga kan se .
alla ytterligare analyser av s�rskilda tekniker , som t.ex. filtersystem , m�ste ta h�nsyn till de tekniska framsteg som skett .
det �r n�dv�ndigt att ge industrin incitament i en s�dan riktning genom internationellt samarbete men ocks� att �ka medvetenheten hos f�r�ldrar , l�rare och barn .
jag vill avsluta med att uppmana medlemsstaterna att forts�tta med den dubbla strategi som f�respr�kats p� gemenskapsniv� , det vill s�ga en strategi f�r " mainstreaming " och s�rskilda �tg�rder till f�rm�n f�r kvinnor .
n�sta punkt p� f�redragningslistan �r debatt om aktuella och br�dskande fr�gor av st�rre vikt .
d�rf�r tror jag att vi om de europeiska institutionerna och europaparlamentet hj�lper det peruanska folket i denna sv�ra situation kan bidra till stabiliteten i landet och bef�standet av de demokratiska institutionerna i hela latinamerika .
herr talman , herr kommission�r ! jag tror det som h�nt i peru visar oss hur l�ngt det ibland kan vara mellan ordens formella betydelse och deras verkliga inneb�rd .
f�r att undvika en katastrof �r det absolut n�dv�ndigt att europa agerar politiskt ocks� p� den sydamerikanska kontinenten .
b5-0789 / 2000 av schroedter med flera f�r gruppen de gr�na / europeiska fria alliansen om situationen i afghanistan .
det verkar som om det helt enkelt handlar om grupper av m�n som befinner sig i en v�rld d�r inget annat r�knas �n deras egen sammanh�llning och deras eget f�rtryck av kvinnorna .
det inneb�r att konflikten �r mycket komplicerad , och att ingen l�sning �r inom synh�ll och �nd� , p� den punkten �r vi eniga , beh�vs det en skyndsam l�sning .
bara en politisk l�sning kan d� g�ra det m�jligt att �terst�lla fred , stabilitet och respekt f�r r�ttigheter .
en del kolleger har redan n�mnt en miljon flyktingar , en miljon invalider till f�ljd av minorna , tusentals kvinnor som �r fr�ntagna sina mest grundl�ggande r�ttigheter , som exempelvis r�tten till utbildning , h�lso- och sjukv�rd , arbete eller r�tten att r�ra sig fritt : det m�ste vara fruktansv�rt f�r m�nga av dessa kvinnor - som var vana vid utbildning , vid en sekulariserad tillvaro - att inskr�nkas p� detta omr�de utan n�gon frihet .
s� l�nge talibanledningen forts�tter att uttala sig tvetydigt betr�ffande kontrollen av opiumplantagerna kommer inte kommissionen att st�dja n�gra drogbek�mpningsprojekt i afghanistan .
men som linkohr tidigare p�pekade , problemet med latinamerika �r just att vi bara �gnar oss �t l�nderna d�r n�r det f�rekommer problem .
sedan dess har situationen blivit �nnu v�rre f�r samh�llena d�r .
b5-0779 / 2000 av dupuis med flera f�r tekniska gruppen f�r oberoende ledam�ter om makedonien .
tyv�rr har det blivit s� att problemet inte f�tt n�gon l�sning p� senare tid under den senaste regeringen fram till 1998 .
det �r en vinst f�r makedonien .
herr talman , mina damer och herrar ! min grupp kommer att st�dja f�religgande f�rslag som vi har undertecknat , f�r jag anser att det �r riktigt att en l�sning som uppn�tts i makedonien och g�r det albanska folket tillm�tes �ven st�ds av europeiska unionen .
av den anledningen har kommissionen vid flera tillf�llen uppmanat makedoniens myndigheter att l�sa den ouppklarade fr�gan om universitetsutbildning p� det albanska spr�ket .
b5-0791 / 2000 av korakas med flera f�r gruppen europeiska enade v�nstern / nordisk gr�n v�nster om fartyget express saminas f�rlisning .
eftersom vi respekterar kammarens beslut i f�rrg�r , har vi g�tt in f�r en kompromiss och vi har kommit fram till en gemensam text , tack vare alla gruppernas uppenbarligen mycket goda samarbetsvilja .
jag skulle vilja s�ga ang�ende resolutionen , eftersom det har framlagts vissa �ndringsf�rslag , att �ndringsf�rslaget om fartygsregister faktiskt �r en punkt som finns med i texten .
under den knivskarpa konkurrens som r�der vid upphandlingar , kan f�retag alltf�r ofta pressas att s�nka kostnaderna , och jag vill inte vara med om att det blir s�kerhetsaspekterna som offras .
det �r desto mer tragiskt eftersom skulden till det �r dispensen fr�n europeiska unionens lagstiftning .
kommissionens uppgift �r att �vervaka den praktiska till�mpningen av dessa r�ttsliga ramar inom ramen f�r sin �vervakningsroll som fastst�lls i f�rdraget .
jag vill p�peka att en m�rklig tendens har uppkommit .
jag vill inte d�lja det faktum att situationen inte �r enkel och att vi kommer att f� uppleva sp�nda �gonblick de n�rmaste dagarna , men vi m�ste alla h�lla huvudet kallt s� att inte situationen �verg�r till en allvarlig konflikt .
segern uppn�ddes trots att regimen gjorde och fortfarande g�r stora anstr�ngningar f�r att f�rhindra den .
vi f�rd�mer � det best�mdaste det �verdrivna och urskillningsl�sa ins�ttandet av v�ld .
i det h�r �gonblicket finner vi att parlamentet i belgrad st�r i ljusan l�ga - vi vet vad det inneb�r att s�tta ett parlament i europas historia i brand , och vi vet ocks� vilket ansvar de ledare har som leder sitt folk i f�rd�rvet .
jag tycket att det var mycket chockerande att se att en ambulansf�rare sk�ts ner vid kravallerna och f�r det andra , d�r jag sj�lv var med , en ambulansf�rare sk�ts i foten fr�n tio centimeters h�ll f�r att han ville hj�lpa m�nniskor .
men �ven den palestinska staten har samma r�ttigheter .
de senaste dagarnas h�ndelser visar emellertid alldeles riktigt p� att fredsprocessen �r synnerligen �mt�lig .
f�r en s�dan situation kr�vs fink�nslighet .
�n en g�ng f�rv�xlar man , � ena sidan , en demokratisk stat som med sv�righet k�mpar mot en mycket sv�r situation med , � andra sidan , auktoriteten mitt i palestina som , f�rvisso inf�r en provokation , anv�nder skjutvapen vid f�rsta b�sta tillf�lle f�r att beskjuta de israeliska ordningsstyrkorna .
kommissionen och r�det kommer att g�ra sitt och det �r det viktigaste som f�r n�rvarande st�r p� dagordningen i jugoslavien ; det har vi alltid varit angel�gna om .
jag vill ocks� s�ga - och det �r egentligen en uppmaning till r�det men jag s�ger det nu till kommissionen och till oss sj�lva - l�t oss inte bara komma med vackra uttalanden om det st�d som vi inom kort vill ge till serbien utan l�t oss ocks� skapa utrymme i v�r egen budget , europeiska unionens budget , s� att vi inom kort inte beh�ver konstatera att vi endast kan hj�lpa serbien genom att ta pengar fr�n andra projekt i balkanomr�det .
s� l�d rapporten kl . 17.53 .
n�r det g�ller f�rh�llandet till unders�kningskommitt�n vill jag ocks� betona att det m�ste vara en internationellt sammanst�lld unders�kningskommitt� och att tydliga gr�nser m�ste l�ggas f�r dess befogenheter .
det skulle vara katastrofalt att helt och h�llet g� �ver till euron under nuvarande omst�ndigheter .
parlamentet skall i dag besluta om en mycket enkel fr�ga , huruvida kroatien skall anslutas till de l�nder som europeiska investeringsbanken kan bevilja l�n som garanteras av eu .
v�r politiska grupp har uppr�tth�llit en strategi i budgetf�rfarandet f�r �r 2001 d�r en klar f�rb�ttring efterstr�vas av kvaliteten p� utgifterna och en f�rb�ttring av kontrollmekanismerna f�r utf�randet .
f�rhoppningsvis skall de hoppfulla signalerna fr�n kroatien och nu �ven fr�n jugoslavien sporra oss att finna en l�sning f�r budgeten och problemen i budgetplanen .
europeiska unionen kan inte till�ta sig att efter de vackra orden i g�r och efter att ha beviljat denna garanti i dag komma till belgrad i morgon med tomma h�nder .
kroatien satte redan f�r tio �r sedan ig�ng med demokratiseringen och med demokratin .
d�rf�r �r det viktigt att kroatien �ntligen f�r ett associeringsavtal som g�r klart att det handlar om ett europeiskt land med blicken entydigt riktad mot anslutning till europeiska unionen .
d�rf�r �r det bra att redan nu s�tta in �tg�rder f�r detta .
i l�mplighetsrapporten om ett stabiliserings- och associeringsavtal med kroatien fr�n maj 2000 kommer kommissionen till slutsatsen att villkoren har uppfyllts f�r att f�rhandlingar skall tas upp med kroatien .
efter m�nga �rs sv�righeter f�r befolkningen - sv�righeter av alla slag - kan vi nu �ntligen p� ett mycket demokratiskt s�tt �ter v�lkomna serbien i folkgemenskapen i europeiska unionen .
finns det n�gra andra synpunkter p� protokollet ?
jag vill att parlamentet skall registrera dessa �vertr�delser och naturligtvis kr�va omval i omr�det kring himara .
fru talman ! det har fallit fler offer f�r eta , men det har ocks� fallit fler offer f�r det spanska f�rtrycket : fler arresteringar , fler torterade , nya utspridningar av politiska f�ngar som f�ngslats i baskien .
jag anser att den minst d�liga l�sningen till sist �r att till�mpa minutregeln , som man f�rresten har kunnat konstatera .
vad g�ller herr le pen , �r det uppr�rande f�r europaparlamentet och alla demokrater att h�ra herr le pen anv�nda ordet " dignitet " .
vi skulle �tminstone �nska att det skulle bli det p� nytt av ett politiskt sk�l .
vad vi nu g�r �r inget annat �n vad vi redan har gjort p� omr�det skog och v�xter , n�mligen att referera till det horisontala direktivet .
och jag citerar ordagrant det brev ni sj�lv , fru talman , l�ste upp i kammaren den 17 maj .
personligen kunde jag inte anm�la detta , eftersom det r�rde sig om partiv�nner som alltid har varit m�ltavlor av politiska sk�l och det d�rf�r skulle verka som om jag talade i egen sak .
vi m�ste kunna se var det g�rs framsteg , dessa m�ste kunna m�tas , och den socialpolitiska dagordningen m�ste f� en central plats i den politiska diskussionen vid det europeiska toppm�tet .
jag �r �vertygad om att europa inte kommer att bli socialt f�rr�n den ekonomiska politiken , konkurrenspolitiken , utrikespolitiken och hela utvidgningsdiskussionen ocks� f�r ett socialt inneh�ll .
jag skulle framf�r allt vilja gratulera fru van lancker , och �ven utskottet f�r syssels�ttning och socialfr�gor och dess ordf�rande till det bet�nkande som vi skall debattera och som �r ett bevis p� europaparlamentets dynamiska och h�ga engagemang f�r den sociala dagordningen .
vi har speciellt f�rbundit oss vid m�let om full syssels�ttning .
jag vill s�ga n�got om arbetstagares r�rlighet .
vi har ocks� kunnat genomdriva n�gra saker p� det sociala omr�det men inte allt , och det h�ngde samman med att amsterdamf�rdraget �nnu inte hade tr�tt i kraft . i det avseendet �r det h�r sociala handlingsprogrammet eller den h�r socialpolitiska dagordningen av mycket stor betydelse .
kommissionen har i sitt meddelande hittat en ram f�r den socialpolitiska dagordningen , som jag tycker anammar andan fr�n toppm�tet i lissabon p� ett bra s�tt .
den br�dskande sociala fr�gan och bevarandet av den europeiska sociala modellen kr�ver initiativ i syfte att inf�ra r�ttigheter till en inkomst , en l�n och hyggliga pensioner f�r alla i europeiska unionen .
jag tror att kraften m�ste komma nedifr�n , och att det g�ller att s�tta in st�det p� den niv� d�r problemen finns .
man har prioriterat byggandet av den gemensamma marknaden : principen om fri r�rlighet f�r tillg�ngar , varor och kapital , inf�randet av regler som styr konkurrensen mellan f�retag liksom statligt st�d .
i bet�nkandet st�r det emellertid litet annorlunda formulerat : eftersom man vid toppm�tet uppmanade till en reformering av den sociala modellen , vill man d�rmed se en f�rst�rkning ; eftersom man vid toppm�tet uppmanar till en befrielse av f�retagen och mer flexibilitet , f�resl�s i bet�nkandet fyra nya eller �ndrade direktiv och en rad lagstiftningsinitiativ .
herr talman , k�ra kolleger ! jag vill s�rskilt lyck�nska tv� av de n�rvarande , f�r det f�rsta v�r kollega anna van lancker till hennes framst�ende bet�nkande , f�r det andra kommission�r anna diamantopoulou till hennes utm�rkta framst�llning .
jag tror ocks� att det �r en stor f�rdel om vi lyckas uppn� att direktivet f�ljs , �ndrat och uppdaterat , som handlar om moderskapsledighet , dvs. att m�drar skall f� hj�lp under graviditeten och ett moderskapsskydd n�r kvinnorna m�ste forts�tta att arbeta under denna tid .
social kvalitet �r inte gratis .
dessa tv� nya politiska inslag genomsyrar hela inneh�llet .
sv�righeten ligger i att den sociala dagordningen , p� grund av f�rdragets r�ttsliga grunder , inte utg�rs av enhetlig lagstiftning eller direktiv med konkreta steg och m�tt f�r medlemsstaterna .
detta arbete har g�tt ganska snabbt , trots att det tog lite tid i b�rjan .
jag s�ger det h�r s� att inte n�gra mystiska , tekniska f�rfaranden g�r att detta missuppfattas .
i enlighet med detta m�ste problemen kring tillg�ngen till social trygghet individualiseras .
den omfattar alla de omr�den p� vilka man beh�ver vidta �tg�rder och , om den samordnas p� ett framg�ngsrikt s�tt , skulle kunna spela en stor roll f�r kvinnor n�r det r�r vardagens alla aspekter .
p� detta omr�de liksom p� m�nga andra �r det absolut n�dv�ndigt att myndigheterna f�rm�r visa en �kta pluralism i valet av sina associerade samtalspartner .
lika tillg�ng till och ett fullst�ndigt �tnjutande av sociala r�ttigheter f�r kvinnor och m�n , vilket skulle inneb�ra att man bevakar till�mpningen av lagstiftningen inom det sociala omr�det i f�rh�llande till mammaledigheter , moderskapsskydd , arbetstider , anst�llningskontrakt , osv .
detta �r en konsekvent till�mpning av gender mainstreaming-konceptet .
herr talman ! jag tycker det vore v�ldigt synd om inte nicole p�ry ocks� tog tillf�llet i akt och uttalade sig nu n�r hon �r h�r , s� att vi kunde f� h�ra hennes synpunkter ocks� .
omr�stningen kommer att �ga rum i morgon kl . 12.30 .
vi f�r helt enkelt se till att �ndra p� detta .
den gemensamma marknaden �r n�dv�ndig n�r det r�r fr�mjandet av konsumenternas intressen .
jag skall ge ett av flera exempel , ett exempel som f�r tillf�llet diskuteras livligt inte enbart i min region .
nu har f�rvisso en del h�nt de h�r dryga 200 �ren , men vi har samma str�vanden idag .
och det �r tydligt att finansministrarna runt om i europa �r mycket mottagliga f�r dessa p�st�enden .
l�t mig avslutningsvis s�ga f�ljande : vi beh�ver en mer exakt definition av den relevanta marknaden , eftersom marknaden alltmer s�llan �r den nationella marknaden .
i forts�ttningen m�ste man komma ih�g att n�r det till exempel g�ller intern konkurrens finns st�d som �r s�rskilt viktiga och v�rdefulla f�r glest befolkade l�nder d�r avst�nden �r l�nga .
i detta sammanhang har ni omarbetat ett meddelande om offentlig service och �nnu en g�ng presenterat det r�ttsliga l�get .
ett hj�rtligt tack g�r till riis-j�rgensen f�r hennes v�rdefulla bidrag i egenskap av f�redragande av den 29 : e rapporten om konkurrenspolitiken .
s�rskilt uppm�rksammade vi den oro parlamentet gav uttryck f�r vad g�ller fr�gorna om �ternationalisering och r�ttss�kerhet .
det vi m�ste arbeta tillsammans f�r , �r att stegvis uppn� en faktisk gemensam marknad p� marknaden , som str�cker sig bortom den nationella marknaden .
jag har allts� endast talat f�r min grupp , inte f�r hela parlamentet .
syftet med denna rapport fr�n kommissionen �r att skapa en grund f�r granskningen av den �vergripande mekanismen f�r medelfristigt ekonomiskt st�d och en eventuell �versyn av denna .
n�sta punkt p� f�redragningslistan �r bet�nkande ( a5-0195 / 2000 ) av kla� f�r utskottet f�r utveckling och samarbete om f�rslag till r�dets direktiv om �ndring av direktiv 68 / 193 / eeg om saluf�ring av vegetativt f�r�kningsmaterial av vinstockar ( kom ( 2000 ) 59 - c5-0090 / 2000 -200 / 0036 ( cns ) ) .
detta inneb�r i klartext att europaparlamentet skulle ge gr�nt ljus f�r experiment med genetiskt modifierade organismer f�r f�r�kning eller f�rb�ttring av vinstockar .
man kan anse att de nya eller aktualiserade best�mmelserna i det f�reslagna direktivet p� ett tillfredsst�llande s�tt uppfyller f�rv�ntningarna hos de yrkesverksamma inom sektorn f�r vinplantskolor och vinodling och att de b�r bidra till en b�ttre kvalitet i de f�reslagna materialen och underl�tta kontrollen av handeln p� marknaden av vinstockar och vinrankor av de organ som har ansvar f�r denna kontroll .
om kommissionen verkar upphetsad �ver kloning och genetisk modifierade organismer f�renade har f�redraganden g�tt �ver i en verklig frenesi och l�gger i begreppet genetiskt modifierade organismer in genotyper som hon finner �verallt .
slutligen kan vi godk�nna �ndringsf�rslag 27 som lavarra och garot lade fram senare .
fru talman ! jag ser under punkt 13 i protokollet " meddelande om f�rverkande av le pens mandat " att ni trodde er kunna uttala er i parlamentets namn , precis som ordf�randen f�r utskottet f�r r�ttsliga fr�gor och den inre marknaden gjort f�r utskottets r�kning .
ni kan kontrollera det i det muntliga protokollet .
n�r det g�ller regeringskonferensen tror jag att arbetet p� ministerniv� f�re biarritz hade kommit s� l�ngt det var m�jligt , och detta informella r�d kom d�rf�r i r�tt tid f�r att bekr�fta vissa framsteg , f�r att ge riktlinjer f�r arbetets slutfas som vi allts� redan har g�tt in i .
de tv� formlerna finns allts� p� bordet , vi m�ste bed�ma dem hur man genom dem kan se till att gemenskapens allm�nna intresse respekteras .
europeiska unionen h�ller fast vid sina �taganden och tog konsekvenserna av denna politiska omv�lvning redan vid r�det ( allm�nna fr�gor ) den 9 oktober , d� man beslutade att h�va sanktionerna , d�ribland oljeembargot och flygembargot , som drabbat f�rbundsrepubliken jugoslavien sedan 1998 , naturligtvis med undantag av sanktionerna som g�ller milosevic sj�lv och hans omgivning . presidenten besvarade allts� ordf�randeskapets inbjudan att komma till biarritz f�r en lunch med stats- och regeringscheferna .
mina damer och herrar parlamentsledam�ter ! n�r det g�ller dessa tv� fr�gor som faktiskt kommer att l�sas f�rst i slutet och f�r vilka vi inte f�r n�gon �verenskommelse alls om vi inte �r �verens om allt , m�ste vi hitta en l�sning .
detta var ett positivt tecken .
r�dets tj�nstg�rande ordf�rande talade om andan i nice .
det �r en viktig fr�ga f�r oss som �r med och f�r dem som kan komma att ansluta sig .
fru talman ! f�r det f�rsta vill jag ber�mma europeiska r�det f�r att det godk�nt f�rslaget till stadga som definitivt .
jag uttrycker ocks� min grupps och en rad icke-statliga organisationers �nskan att f� se stadgan utvecklas , forts�tta att f�rb�ttras , bl.a. f�r att garantera skydd av r�ttigheterna och mer effektiva r�ttigheter f�r unionens medborgare , f�r de anst�llda , f�r medborgare i tredje land och f�r de utslagna .
det handlar om det enda s�ttet att �teruppr�tta en verklig balans med de olika institutionerna i v�r europeiska union .
man kunde ha hoppats p� lite vackrare v�der , men jag tror att det var lite b�ttre �n vad kommission�ren sade inom europeiska r�det , som jag deltog ifr�n b�rjan till slut .
det handlar verkligen om att f�rst�rka gemenskapsramen .
det �r den f�rsta texten fr�n europeiska unionen som medborgarna kan konsultera utan att k�nna sig fullst�ndigt fr�mmande inf�r dess inneh�ll .
jag anser hur som helst , fru talman , att m�tet i biarritz har tillf�rt n�got mycket positivt : ett enh�lligt godk�nnande av stadgan .
det �r anledningen till att man talar s� mycket om sm� och stora stater .
men vi m�ste snarast f�rse unionen med denna stadga .
d�rf�r f�rhandlade man a minima . vi har en minimal stadga , s�rskilt n�r det g�ller de sociala r�ttigheterna .
vi vet alla att utvidgningen av unionen inte kan �ga rum f�rr�n beslutsprocesserna inom de stora institutionerna har �ndrats . en s�dan reformprocess m�ste dock vara r�ttvis och balanserad .
v�r debatt i dag har f�rresten samma st�mning .
man kan ocks� notera framsteg i fr�ga om artikel 7 , om hur man skall agera , d� europeiska unionens grundl�ggande v�rden kr�nks .
en annan fr�ga g�ller kommissionens reformering .
de stora l�ndernas krav p� �kad makt i r�det och parlamentet skulle , om de tillgodos�gs , rubba hela balansen inom eu och inneb�ra att de sm� l�nderna fick betala hela priset f�r utvidgningen .
den tragiska utvecklingen i mellan�stern har naturligtvis gett upphov till ett oerh�rt bakslag , och de senaste dagarnas v�ld , det stora antalet offer , har naturligtvis v�ckt starka k�nslor i den allm�nna opinionen i europa och h�r i parlamentet . och med r�tta .
herr talman , �rade kolleger ! det �r synd att bar�n crespo inte �r n�rvarande i kammaren efter at ha sagt vissa saker om den politiska kraft som jag f�retr�der .
men vi b�r ocks� titta p� v�r egen situation .
vi m�ste inse att de sm� staterna i en statsunion �r j�mst�llda med de stora staterna , och att vi m�ste kompensera de stora staterna p� annat s�tt .
jag har f�rst�tt att handlingen har tagits emot v�l i biarritz , och att den efter n�gra juridiska f�rtydliganden kan godk�nnas via ett officiellt uttalande av toppm�tet i nice f�r att i framtiden bli upptagen i f�rdragen .
fr�gan �r d�remot om alla l�nder f�r en kommission�r samtidigt , och om vi d�rmed f�r en stor - och en dag en mycket stor - kommission , som naturligtvis m�ste omorganiseras , eller om det blir " inte alla p� en g�ng " .
jag n�mnde nyss mycket exakt n�gra av de best�ndsdelar som kommer att g�ra det m�jligt f�r oss att omedelbart inse om reformen �r tillr�cklig eller otillr�cklig .
muntlig fr�ga till kommission ( b5-0543 / 2000 ) i enlighet med artikel 42 i arbetsordningen fr�n napolitano f�r utskottet f�r konstitutionella fr�gor om artikel 158 i eg-f�rdraget om �ars st�llning .
n�r freden v�l garanterats b�rjade �steuropa att sk�ta sina �taganden genom att str�va efter v�lst�nd .
vi vill ha en verklig konstitution .
jag har haft gl�djen , herr talman , att konstatera att de f�rslag som p� senare tid har lagts fram till regeringskonferensen i huvudsak sammanfaller med alla eller en del av de krav som jag har tagit upp . jag hoppas att anden i biarritz - som �beropas i dag - materialiseras , f�r de andar som inte materialiseras f�rvandlas till sp�ken och det vimlar av s�dana sp�ken p� loftet till den europeiska byggnaden .
vi beg�r inget konkret och framf�r allt , vi beg�r inga bidrag : vi beg�r att denna princip om �karakt�ren skall erk�nnas av alla , s� att unionens medborgare har samma f�ruts�ttningar fr�n b�rjan , s� att alla skall f� samma m�jligheter att n� �nda fram .
man kan d�rf�r knappast s�ga att allt fungerar exakt som om vi var femton , jag ber om urs�kt f�r att jag betonar en s�dan sj�lvklarhet .
jag tror att vi verkligen kan tala om en konstitution , och planera f�r villkoren f�r hur den skall skrivas , f�rst n�r vi vet vad vi vill placera i den .
flera av er , men �ven medlemsstaternas representanter , har redan sagt att den traditionella formuleringen fr�n regeringskonferensen sannolikt inte var den b�sta .
n�r det g�ller den id� ni tog upp att introducera denna debatt i regeringskonferensen , f�refaller det mig uppriktigt sagt , herr segni , med tanke p� omfattningen och sv�righeten med de �vriga fr�gorna som st�r p� dagordningen f�r denna regeringskonferens , att det skulle vara mer l�mpligt att , s�som gjorts tidigare f�r andra materiella felaktigheter i artiklarna i f�rdragen , komma fram till en r�ttelse av texten enligt f�rfarandet i wienkonventionen om f�rdragsr�tten , f�r att konkret och precist j�mf�ra de olika spr�kliga versionerna av denna artikel .
efter�t kommer det inte l�ngre att finnas n�gra krav fr�n v�r sida .
� andra sidan f�r det inte utg�ra ett hinder f�r utbytet eller �stadkomma en uppdelning av den gemensamma marknaden , ett avbrott i solidariteten och sammanh�llningen mellan medlemsstaterna , eller s�som kommission�r barnier sade , en s�nderdelning av gemenskapens regelverk .
efter nice-m�tet , som vi alla hoppas blir framg�ngsrikt , �r det viktigt att ta detta n�sta steg f�r att skapa en mer demokratisk union .
nu skall jag g�ra vad jag kan f�r att �vertala mina landsm�n att f�ra denna stafettpinne vidare under sveriges ordf�randeskap .
det f�r n�mligen inte vara s� att bara de femton medlemsstaterna diskuterar och beslutar om en f�rfattning , n�r vi ju alla vet att vi i slutet av detta �rtionde kommer att ha ett europa med 27 medlemsl�nder !
men om det �r tillsammans �r det n�dv�ndigtvis samtidigt .
argumentet mot detta och varningen f�r ett europa med flera hastigheter kommer jag fortfarande ih�g .
f�r det f�rsta ang�ende metoden , ett f�r allm�nheten utt�mt f�rfarande som faktiskt �sidos�tter unionens �vriga institutioner och d�r regeringarna blivit offer f�r sin egen labyrint .
herr talman ! vi har h�rt att man har gjort framsteg i biarritz om �kat samarbete .
� andra sidan finns det en risk f�r att det n�rmare samarbetet fr�n ett annat h�ll kommer att uppl�sa europas enhet och leda oss till en hel mosaik av olika samarbetsformer mellan regeringar .
jag medger dock att de politiska f�ruts�ttningarna inte har funnits f�r att g� l�ngre , och d�rf�r godk�nner jag utan reservationer duhamels bet�nkande som vi nu debatterar .
som sista talare skulle jag vilja gratulera b�de duhamel till hans utomordentliga arbete och gil-robles till hans eget arbete .
d�rf�r vill vi ha �rendet �terf�rvisat till oss .
det tar jag inte h�nsyn till .
vad inneb�r uttrycket " den tidsperiod inom vilken medlemsstater skall garantera arbetsl�sa tillg�ng till syssels�ttningspolitiska �tg�rder inte b�r �verstiga tv� �r " , om inte ett hot mot arbetsl�shetsunderst�det ?
herr talman ! jag r�stade f�r souchetbet�nkandet som syftar till att i st�rre omfattning till�ta att man f�rvandlar jordbruksprodukter till f�rpackade livsmedel .
varf�r ? d�rf�r att bet�nkandet godk�nner m�jligheten att g�ra om vinstockar till genetiskt modifierade organismer och d�rmed , i morgon , till�ter att vi dricker genetiskt modifierat vin .
enligt ett f�rslag skall man till�ta saluf�ring av f�r�kningsmaterial f�r vinstockar med l�gre s�kerhetskrav , n�r det uppst�r tillf�lliga sv�righeter , men man definierar inte vilka sv�righeter det i s� fall skulle r�ra sig om .
sk�let �r att mr . smith betalar litet i pensionsavgift , medan det som signor rossi betalar �r mycket mer .
i princip kan en decentraliserad till�mpning av gemenskapslagstiftningen bara bli framg�ngsrik om det finns starka fasta �taganden om att detta kommer att till�mpas enhetligt �ver alla europeiska unionens territorier .
statliga st�d har traditionellt anv�nts av medlemsstater som instrument f�r industri- och socialpolitik .
jag �r inte lika n�jd med den tanke som omn�mns i punkt 2 om att det statliga st�det inte f�r stiga .
jag anser det oacceptabelt med de p�tryckningar och andra liknande �tg�rder som f�resl�s , t.ex. om registrering och utv�rdering av " effekterna " av de statliga st�d�tg�rderna .
avsnitt v , revisionsr�tten
till och med kommissionen har varit mycket �terh�llsam n�r det g�ller att f�resl� betalningar i f�rslaget till budget , alltf�r �terh�llsam anser vi .
detta m�ste motverkas p� alla politiska niv�er , lokalt , regionalt , nationellt , men ocks� europeiskt .
efter den gl�djande utg�ngen av valen i serbien skall vi nu ocks� st�dja serbien med finansiella medel och inte bara med vackra ord i s�ndagspredikningar .
f�r det tredje : skattebetalarnas pengar m�ste i slut�ndan ge ett merv�rde .
vi �r ju direkt bundna till europeiska centralbankens r�ntesats , och vi f�resl�r d�rf�r att man forts�tter p� den inslagna politiken i fr�ga om byggnaderna , eftersom detta bidrar till att snarast m�jligt befria oss fr�n dessa r�nteb�rdor .
ett stort sorgebarn �r fortfarande ekonomiska och sociala kommitt�n .
herr talman , mina damer och herrar ! i juni 2002 l�per eksg-f�rdraget ut .
det tycks oss vara absurt , eftersom det fortfarande kommer att finnas en driftsbudget under andra halv�ret 2002 , och vi vill d�rf�r ha en granskning av f�rh�llandet mellan omplaceringsst�den och det sociala bist�ndet .
det f�rslag jag ber er godk�nna , genom att r�sta f�r bet�nkandet , utg�r kulmen p� en l�ng process och svarar mot en ur�ldrig str�van hos parlamentet .
vi anser att detta uttalande b�r ing� i det interinstitutionella avtalet , men hur som helst vill jag p�peka f�r er att det endast �r meningsfullt inom ramarna f�r ett interinstitutionellt avtal som har en budgetplan .
jag hoppas att budgetarbetet genomf�rs i samma anda , s� att vi kan uppn� en budget , f�r budget�ret 2001 , som ger oss m�jlighet att m�ta de prioriteringar och utmaningar som v�ntar europeiska unionen inom kort .
n�r det g�ller besparingen p� 225 miljoner euro inom landsbygdsutveckling tas det i r�dets st�ndpunkt h�nsyn till de f�rseningar som ackumulerats i de nationella utvecklingsplanerna f�r landsbygden .
jag antar att det ocks� �r �verdrivet .
det vi beg�r av medlemsstaterna g�ller ocks� f�r den europeiska budgeten , och att komma �verens om allt detta g�r budgetpolitiken s� sp�nnande , vilket alla vet som �gnar sig �t den .
det har bland annat formulerats villkoret att kommitt�f�rfarandet skall �ndras .
fr�gan om man kan lyfta ut de n�dv�ndiga �tg�rderna ur det hittillsvarande f�rslaget f�r programmet f�r medelhavsomr�det �r en politisk och inte n�gon teknisk fr�ga .
vi skall st�dja hans och chris pattens f�rs�k att st�rka kommissionens handlingskraft genom parlamentets kunskaper och genom den n�dv�ndiga parlamentariska kontrollen , som ju inte g�ller r�det och solana .
den f�rsta g�ller genomf�randet av ett pilotprojekt avsett att finansiera en informationskampanj inom de femton medlemsstaterna mot den brottsliga pedofilfarsoten .
h�r har utskottet f�r ekonomi och valutafr�gor st�llt kravet p� ett expertutl�tande f�r att f� l�mplig r�dgivning fr�n europeiska centralbanken i penningfr�gan .
de f�rslag som lagts fram av v�rt utskott och som st�tts av budgetutskottet �r mycket b�ttre .
den som p�st�r att det kanske handlar om att f�rhindra fusioner eller stoppa globaliseringen , s�ger detta enbart av polemiska sk�l .
det �r denna kammares ansvar att st�dja dessa fr�gor i omr�stningen denna vecka , att visa dess fortsatta �tagande f�r att skydda milj�n ock f�rb�ttra folkh�lsan .
fiskeriutskottet som med kommissionen delar principen om budgetstringens , har accepterat de gr�nser som denna anger i sitt prelimin�ra f�rslag och har framf�rt sin oro betr�ffande vissa budgetposter .
att var och en �tar sig sitt ansvar och uppfyller sin skyldighet .
europeiska kommissionen har knappt kunnat klara av utvidgningen av prioriteringarna , och detta har lett till oacceptabla eftersl�pningar vid genomf�randet av �tagandena som g�rs under trycket fr�n allt st�rre budgetar f�r st�d till utl�ndska hj�lp- och samarbetsoperationer .
vi b�r ocks� ha i �tanke att allt detta h�r samman med den kamp mot v�ld i hemmet som bedrivs genom programmet daphne .
det finns inga b�ttre bevakare av f�rdragen �n de europeiska medborgarna .
ramen f�r v�r debatt i dag �r att vi m�ste anv�nda varje m�jlighet vi har i v�r budget f�r att se till att v�ra europeiska institutioner �r redo f�r n�sta etapp av utvidgningen , s�v�l vad g�ller institutionernas strukturer som ett b�ttre s�tt att bedriva politik .
innan jag kommer till det , ett ord om de brittiska konservativas st�ndpunkt .
vi f�rst�r att det finns ett behov av mer personal , men det som �r mest angel�get f�r oss �r att inte bevilja denna beg�ran f�rr�n reformen av institutionerna �r ordentligt i g�ng .
men hit h�r ocks� att man naturligtvis ocks� h�r i m�nga fall skall ge skattebetalaren klart besked , s� att han f�r en faktisk bild av vilka villkor vi arbetar under .
men vi har gamla l�ften respektive tillk�nnagivanden , gemensamt formulerad politik , som senare n�gon g�ng ocks� faktiskt m�ste inl�sas i form av betalningar .
jag vill tydligt s�ga att jag anser att det �r ansvarsl�st om vi ger de m�nniskor som drabbas av katastrofer det intrycket att vi d�rmed skulle kunna l�sa alla problem som h�nger samman med katastroferna .
�ven om vi inst�mmer i kritiken mot r�det p� flera punkter , kan det konstateras att denna strategi skulle inneb�ra en konfrontation d�r ingen f�rlikning �r m�jlig , och som skulle undergr�va de europeiska institutionernas trov�rdighet .
vi befarar att utskottsmajoriteten genom taktik har l�st sig .
haug , v�r huvudf�redragande , f�rs�kte ocks� hon i g�r kv�ll att �ndra sitt bet�nkande p� denna punkt f�r att bem�ta den oro som uttrycktes av min grupp . det tackar jag henne f�r .
avsev�rda besparingar �r m�jliga , vare sig de beror p� att vissa program underutnyttjats eller p� att europeiska unionen �ntligen valt att sluta anv�nda budgetposterna f�r europapropaganda .
vi m�ste ge kommissionen chansen att genom ut�kning av personalen arbeta bort eftersl�pningen .
skatteb�rdan m�ste d�rf�r s�nkas procentuellt , och h�gre statsint�kter kan bara uppn�s via ett ekonomiskt uppsving och den d�rmed f�rknippade ekonomiska tillv�xten .
behoven �r uppenbara , �tagandena �r m�nga , det externa samarbetet f�r att h�vda europeiska unionen �r tydligt , men genomf�randet av flera program �r mycket l�gt .
vi f�rs�ker s�kra parlamentets prioriteringar i utgiftsomr�de 4 .
vi anser att vi har mer vetenskapliga bevis �n er gissning om en siffra .
( skratt och appl�der )
det f�r exempelvis inte vara s� att " de sm� l�nderna " , ett fullst�ndigt opassande uttryck , tror att de kommer att uteslutas fr�n det n�rmare samarbetet , att det n�rmare samarbetet skall betyda f�rtrupp , gravitationscentrum , pionj�rgrupp och att den kommer att vara sluten .
jag tror d�rf�r att det var fullst�ndigt relevant att i detta sammanhang be en extern myndighet som �r moraliskt of�rvitlig att vidta dessa �tg�rder .
n�r det g�ller de konkreta m�jligheterna f�r den colombianska regeringen att undanr�ja de paramilit�ra grupperna �ligger det de colombianska myndigheterna att fastst�lla dem .
m�nga anser att problemen i colombia , liksom i andra l�nder i latinamerika , bottnar i b�ndernas �gande eller icke-�gande av marken .
. ( fr ) jag tror att jag just besvarat fr�gan .
jag vill inte att ni skall tro att r�det inte besvarar de fr�gor det f�r .
kan r�dets ordf�randeskap ange , mot bakgrund av de diskussioner som r�det kan ha haft med ekonomi- och finansministrarna i unionens medlemsstater liksom i tredje l�nder , var motst�ndet mot denna skatt kommer ifr�n och vilka som , enligt r�dets f�rmenande , �r de huvudsakliga politiska och tekniska hindren f�r att det skall kunna inf�ras en s�dan skatt ?
inr�ttandet av en tobin-skatt �r frestande . den f�rsvaras p� m�nga h�ll , till v�nster och h�ger , av olika organisationer , politiska eller andra , av icke-statliga organisationer , av universitetsgrupper .
herr ordf�rande !
jag beklagar .
d�rf�r kan de ibland inte urskilja den som �r r�dets tj�nstg�rande ordf�rande .
n�r allt kommer omkring �r fr�gan som jag , personligen , st�ller mig , just h�r , med min impuls som militant , vad som kr�vs f�r att det skall fungera .
r�det forts�tter aktivt granskningen av kommissionens f�rslag samt de n�mnda �ndringsf�rslagen , i syfte att mycket snabbt kunna utarbeta en st�ndpunkt i �rendet .
. ( fr ) jag hoppas att parlamentsledamoten inte blir arg p� mig f�r att jag inte i detalj vill inleda en debatt om bse , som verkligen vore p� sin plats h�r i kammaren , efter att ha haft en debatt om tobin-skatten .
tack f�r ert svar , herr ordf�rande , men fr�gan gick l�ngre �n s� .
herr talman , fru kommission�r ! jag skulle vilja b�rja med att framf�ra mina komplimanger till f�redraganden .
d� k�nde man inte till att r�det och kommissionen av dessa pengar lovar st�d f�r �teruppbyggandet av serbien och kosovo .
det finns fattiga i europa , om det s� bara g�ller pensionerade lantbrukare .
de externa behoven avsl�jar knappheten i kategori 4 .
vi befinner oss nu i f�rsta behandlingen och ni har gott om tid att s�ka uppn� ett fullst�ndigt samf�rst�nd med parlamentet .
vi kan bara vara �ppna och redovisningsskyldiga om alla beslutsfattare �r tydliga om budgeten och besluten bakom budgeten .
som folkvald gl�der man sig naturligtvis �ver varje �tg�rd som kan g�ra budgeten mera begriplig .
d�remot finns det ett folkligt krav p� att vi skall finna en l�sning och st�dja serbien .
jag v�lkomnar tillf�llet att ge ett kort bidrag till denna viktiga debatt och att tala om vikten av jordbruksbudgeten och dess betydelse f�r inte bara b�nder utan f�r samh�llet i stort .
herr talman , kolleger , fru kommission�r ! f�rst och fr�mst vill jag naturligtvis tacka alla f�redragandena .
herr talman ! med sitt budgetf�rslag f�r 2001 har r�det verkligen �vertr�ffat sig sj�lvt .
den politiska stabiliteten h�nger ihop med om levnadsvillkoren kommer att f�rb�ttras .
med tanke p� att kommissionen sj�lv har medgett att medlemsstaternas beg�ran f�r 2001 om betalningar till strukturfonderna �verstiger ber�kningarna i det prelimin�ra budgetf�rslaget med 8 000 euro , tror jag att det nu �r dags att r�det p� fullaste allvar b�rjar �verv�ga att g�ra n�got �t betalningarna och inte �ka de utest�ende �tagandena .
innan denna punkt har klarlagts och diskuterats ing�ende , v�grar jag helt enkelt att �verhuvud taget tala om n�gon revidering av budgetplanen .
finansministrarna fick ju tillbaka betydligt st�rre summor ur fjol�rets budget .
f�r sverige skulle detta medf�ra cirka 65 miljoner euro .
v�r grupp riktar strategin f�r den allm�nna budgeten mot utgifternas kvalitet och effektivitet i budgetstyrningen . det g�ller �ven eksg : s budget .
men min huvudpunkt g�ller avs .
snarare m�ste dessa st�d minskas stegvis . detta under f�ruts�ttning att de ber�rda jordbrukarna garanteras strukturbidrag f�r att st�lla om sin produktion .
jag s�ger utan urs�kt att jag skall ta upp de effekter som europeiska unionen har gett i min region .
den europeiska modellen betraktar skydd av personuppgifter som en grundl�ggande r�ttighet , garanterad av normer som har rang av lag , inspirerade av principen om sj�lvbest�mmande n�r det g�ller information , dvs. den princip enligt vilken var och en skall sj�lv kunna best�mma om och hur de data som r�r vederb�rande f�r samlas in och anv�ndas .
jag litar p� att det t�lmodiga arbete som genomf�rts skall f� fullt st�d av parlamentet och av r�det .
jag hoppas verkligen att man ser till att best�mmelserna inte kommer att till�mpas p� detta s�tt .
enligt min uppfattning �r det klart att det skulle inneb�ra att man d�ljer ansiktet om man skapar en s�dan myndighet enbart f�r gemenskapsomr�det , medan de huvudsakliga problemen , �ven i framtiden , ocks� kommer fr�n organisationer inom den tredje pelaren .
det verkar som om f�redraganden gjort allt som g�r f�r att , framf�r allt i framtiden , ut�ka m�jligheterna att �tminstone samarbeta och eventuellt ocks� p�verka denna fr�ga , varf�r vi ger v�rt fulla st�d till detta bet�nkande .
n�r det g�ller mer specifikt �ndringsf�rslagen i paciottis bet�nkande �r kommissionens st�ndpunkt f�ljande .
den europeiske tillsynsmannen kommer att spela en mycket viktig roll n�r det g�ller gemenskapsinstitutionernas respekt f�r best�mmelser som skyddar medborgarnas personuppgifter .
azorerna , kanarie�arna , guadeloupe , guyana , madeira , martinique och r�union utg�r en speciell enhet vars odelbarhet erk�nns i amsterdamf�rdraget p� grundval av ett nyskapande koncept , de yttersta randomr�dena .
f�r att den nya gemenskapsstrategin till f�rm�n f�r unionens yttersta randomr�den skall fungera kr�vs �tg�rder med inriktning p� de strategiska omr�dena i v�rldskonkurrensen : transport , energi , milj� , informationssamh�llet , forskning eller teknisk utveckling .
vi hoppas att kommissionen kommer att utveckla denna kalender eller detta program och vi hoppas framf�r allt att den stora institution som kommissionen f�r n�rvarande har , den enhets�verskridande gruppen , uppr�tth�ller kontakten med de yttersta randomr�dena och informerar de centrala myndigheterna om v�ra s�rskilda behov och problem .
faktum �r att det vi s�ger i dag och r�star fram i morgon kommer att skapa rubriker i pressen i de sju yttersta randomr�dena och de regionala tv-kanalernas nyhetss�ndningar kommer att informera utf�rligt om det vi s�ger och beslutar h�r .
d�rf�r �r det sv�rt f�r oss att skapa rikedom och syssels�ttning .
jag gl�ds d�rf�r �t att utskottet f�r regionalpolitik visat prov p� dj�rvhet och ambition n�r det g�ller det statliga st�det , beskattningen och konsekvenserna med anledning av utvidgningen .
p� grund av permanenta , of�rdelaktiga omst�ndigheter �r de yttersta randomr�denas s�rst�llning och exceptionella st�d befogat , men man b�r �nd� inte j�mna ut skillnaderna med best�ende begr�nsningar av regler f�r den inre marknaden eller konstant f�retr�de till de strukturella fonderna .
herr talman ! detta parlament - och s�rskilt utskottet f�r regionalpolitik , transport och turism - har varit den stora p�drivaren f�r att anta s�rskilda politiska strategier och program f�r gemenskapens yttersta randomr�den .
det g�r att de kr�ver en s�rskild behandling som tar sig uttryck i en varaktig vilja i en rad �tg�rder .
de l�mnade d�rf�r sitt fulla st�d , i samband med f�rberedelserna av den f�reg�ende regeringskonferensen , till f�rhandlingarna som ledde till att artikel 299.2 antogs - jag har ett mycket exakt minne av det , eftersom jag d� var frankrikes f�rhandlare f�r amsterdamf�rdraget .
vi m�ste f�r �vrigt i sinom tid g�ra samma anstr�ngningar i form av st�d och signaler n�r det g�ller r�det .
herr pohjamo ! nyss tog ni sj�lv upp denna oro genom att h�nvisa till sanchez arbete och engagemang och jag ber er framf�ra v�ra h�lsningar om god b�ttring , med tanke p� hans h�lsoproblem f�r n�rvarande .
en partnerskapsdag h�lls den 23 november 1999 med ett stort antal deltagare .
jag vill inte ta upp den fr�gan p� nytt .
herr talman ! kollegan evans �terkom just till omr�stningen i g�r f�rmiddag , framf�r allt den omr�stning d�r vissa �ndringsf�rslag godk�ndes med en marginal p� bara en r�st .
vi �r vad vi �ter - och sorgligt nog st�mmer det i mitt fall .
det �r fallet med det f�retag som tillverkade poliovaccin i f�renade kungariket med ett serum fr�n kalvfoster , vilket �r f�rbjudet sedan 1999 , och med distributionen av tusen kilo k�tt fr�n bse-smittade djur i en fransk kedja f�r livsmedelsdistribution .
beslutsprocessen m�ste vara klar och �ppen .
herr talman ! f�rst vill jag varmt gratulera f�redraganden bowis , men �ven s�ga till kommission�r david byrne att vi uppskattar det arbete han har f�reslagit oss med denna vitbok samt de f�rbindelser som han uppr�tth�ller med parlamentet , i syfte att f�r framtiden f�rbereda b�sta m�jliga lagstiftning p� omr�det f�r livsmedelss�kerhet .
den dagen kommer vi inte att k�nna n�gon s�rskild stolthet �ver v�ra tidigare rutiner .
dessa �tg�rder �r intimt sammanl�nkade med livsmedelsmyndighetens kommande verksamhet .
i bet�nkandet g�rs mycket riktigt �tskillnad mellan � ena sidan riskbed�mning och � andra sidan riskhantering .
likafullt , herr talman , l�t mig betona en eller tv� punkter .
vem kan slutligen b�ttre �n staterna informera befolkningen om vilka risker som h�nger samman med olika produkter ?
who t�cker hela europa men har d�rut�ver ett vidare ansvarsomr�de som str�cker sig �ver hela planeten , vilket �r viktigt .
det �r f�rnuftigt , s� att den europeiska livsmedelsmyndigheten ocks� kan verka oberoende av kommissionen och d�rigenom - om det skulle kr�vas - hantera kriser s� snabbt som m�jligt .
jag har lagt fram ett f�rslag i den fr�gan och ber er st�dja det f�rslaget .
det som d�r beh�vs �r inte s� mycket vi och kommissionen utan d�r beh�vs medlemsstaterna , f�r de har inte sk�tt sina uppgifter hittills .
min grupp st�der de flesta �ndringsf�rslagen .
ett tydligt regelverk , definitionen av godtagbara risker och ett konkret v�rnande om m�ngfalden livsmedel och lokal produktion �r aspekter som �terst�r att bena ut , liksom skyddet f�r sm� och medelstora f�retag och utbildning av deras anst�llda .
hade en dioxinkris eller en bse-kris kunnat f�rhindras med en europeisk livsmedelsmyndighet ?
det finns ett ouppl�sligt samband mellan att �ta sunt och att �ta gott , ett samband som konsumenterna m�ste g�ras �n mer medvetna om . vi m�ste fr�mja kvalitet och st�dja de typiska lokala produkter som �r en stor rikedom f�r de europeiska folken .
d�rf�r kommer vi ocks� - som min kollega mihail papayannakis sade - att godk�nna och st�dja bet�nkandet .
dessutom b�r inga livsmedel som har modifierats genetiskt eller inneh�ller genetiskt modifierade ingredienser till�tas i livsmedelskedjan f�rr�n de har testats ordentligt , och d� endast med tydligt angiven m�rkning .
kolleger , herr talman ! i och med den h�r vitboken om livsmedelss�kerhet har en viktig grund lagts f�r b�ttre mat i framtiden och �ven f�r en milj�- och m�nniskov�nligare livsmedelsproduktion , hoppas jag .
f�r att konsumenternas tillit till att livsmedlen �r s�kra skall kunna �teruppr�ttas och bibeh�llas m�ste livsmedelsmyndigheten inleda sin verksamhet med tillr�ckliga offentliga resurser .
herr talman ! jag vill gratulera john bowis till ett gott arbete .
sj�lv t�nker jag inte s� , utan jag litar p� den europeiska integrationsid�ns kraft och grundprinciper inom hela eu-omr�det .
dessutom kommer en del av myndighetens �ndam�lsenlighet att ligga i en �ppen beslutsprocess och snabba offentligg�randen p� internet av dess unders�kningsresultat och yttranden , i likhet med till exempel det f�rtr�ffligt v�l fungerande food and veterinary office i dublin .
jag v�lkomnar det f�rh�llandet att det r�der en bred enighet om huvudprinciperna : att ett nytt vetenskapligt organ med ansvar f�r riskbed�mning i fr�ga om livsmedelss�kerhet b�r inr�ttas , att det skall vara oberoende , ansvarsskyldigt , erbjuda insyn och omfattas av de krav objektiv forskning och aff�rsm�ssig sekretess st�ller , och att det b�r f�rse allm�nheten med l�ttillg�nglig och begriplig information .
allas erfarenheter och kunskaper kan samlas h�r och kunskaperna kan utnyttjas i hela europa .
vi har vetenskapliga kommitt�er som ger r�d �t kommissionen .
redan betr�ffande huvudfr�gan i vitboken , inr�ttandet av en myndighet f�r livsmedelss�kerhet , r�der h�gst motstridiga uppfattningar .
det prioriterade och absoluta intresset f�r m�nniskan grundar sig p� dessa principer .
efter att den godk�nts i medlemsstaterna och h�r i parlamentet skall vitboken ocks� f� en lagstiftande form i ett nytt f�rslag till direktiv .
flera f�rslag har redan lagts fram f�r r�det och parlamentet , exempelvis paketet med f�rslag om en omarbetning och uppdatering av lagstiftningen om hygien .
jag finner det uppmuntrande att se den h�ga graden av samst�mmighet mellan parlamentets synpunkter , s�som de formuleras i det f�rslag till bet�nkande som ni nyss har diskuterat , och sj�lva vitboken .
. ( it ) herr talman , herr kommission�r , ledam�ter ! det �r inte f�rsta g�ngen detta parlament �gnar sig �t fr�gan om landminor .
den sista punkten g�ller �ndringsf�rslagen .
d�rf�r m�ste vi beklaga det faktum att en medlemsstat , finland , inte har undertecknat den , och att en annan , grekland , �nnu inte har ratificerat den , vilket v�r kollega luisa morgantini precis har n�mnt .
utmaningen �r enorm , men omf�nget av detta drama kr�ver en anstr�ngning och ett enormt arbete f�r att f� slut p� situationen .
n�r allt kommer omkring var det europaparlamentet som gick i spetsen f�r unionens kamp mot truppminor .
europeiska unionens st�ndpunkt �r tydlig och lades fast i 1997 �rs gemensamma �tg�rd f�r att bredda anslutningen till och ratificeringen av ottawakonventionen till att omfatta s� m�nga l�nder som m�jligt .
vi har antagit en strategi som �r flexibel och samordnande snarare �n rigid och centralstyrd .
p� samma s�tt vill vi inte skapa n�gon ny kommitt� , om det s� vore en f�rvaltningskommitt� eller en r�dgivande kommitt� .
regeringar har gjort utf�stelser och utlovat stora summor pengar .
kommission�ren med ansvar f�r yttre f�rbindelser har tidigare erk�nt att kommissionens yttre bist�ndsprogram har varit ett bekymmer .
herr kommission�r ! ni s�ger : jag �r emot ett antal �ndringsf�rslag .
bonino och patten har r�tt i att det �r sj�lvklart att man skall f�rst�ra lagren , eftersom det bara kostar en hundradel att f�rst�ra en lagrad mina i j�mf�relse med vad det kostar att f�rst�ra en mina som �r utplacerad p� ett st�lle d�r man har sv�rt att hitta den .
eu : s alla organ m�ste agera initiativkraftigt och p� s� s�tt att de fattiga l�nder som lider mest av minproblemet effektivt f�s med i programmet .
att undanr�ja minor �r inte l�ngre ett milit�rt problem , utan en ytterst viktig humanit�r fr�ga .
jag vill uttryckligen po�ngtera att det �r n�dv�ndigt att uppmana ytterligare stater att ansluta sig till ottawakonventionen och i vissa fall snabbt ratificera denna f�r att m�jligg�ra en internationell samordning liksom en rehabilitering av offren .
d�rf�r yrkar jag p� att r�det , som inte �r n�rvarande h�r , och kommissionen , meddelas hur betydelsefullt det �r att beloppet �kas , med tanke p� att f�r varje mina som elimineras placeras tyv�rr mellan 20 och 50 nya ut .
vi f�r inte f�r den skulle gl�mma bort att europeiska unionen , och i synnerhet europaparlamentet , har �nnu b�ttre m�jligheter att unders�ka vart v�ra finansmedel p� det omr�det egentligen tar v�gen .
m�nga av offren �r sm� barn , fruktansv�rda intryck , hemska stympningar som f�rst�r deras levnadsbana innan de knappt har hunnit p�b�rja denna .
jag skulle � min sida s�rskilt vilja betona att f�rdraget b�r generaliseras �nda tills det blir en fullst�ndig framg�ng , f�rst och fr�mst genom att de olika staternas lagar skall bringas i �verensst�mmelse med f�rdraget , s� att vi inte f�r ett nytt exempel p� ett internationellt avtal som inte kommer att till�mpas .
kritiken inneh�ller dock skenhelighet och okunskap .
detta arbete m�ste ocks� bli effektivare genom samordning och kontroll av processerna och genom att ge de icke-statliga organisationerna en st�rre roll .
i bet�nkandena trycker man mindre p� det faktum att de flesta minor har tillverkats i andra l�nder �n d�r de gr�vs ned .
jag kan bara f�rfasa mig om kommissionen verkligen g�r in f�r att st�dja dessa nyss godk�nda , helt orealistiska , i det n�rmaste absurda krav .
kommissionen kommer att utnyttja sin intiativr�tt och st�dja medlemsstaterna f�r att f� till st�nd n�dv�ndiga f�r�ndringar .
flera av kraven i van lanckers bet�nkande �r inte godtagbara .
bakom de juridiska h�rklyverierna fr�n olika h�ll och kanter bekr�ftade toppm�tet i biarritz att europas utvidgning best�r av en besv�rlig kohandel .
- ( de ) vi i frihetspartiet har redan fr�n b�rjan uttalat oss f�r en stadga f�r de grundl�ggande r�ttigheterna och f�r att denna skall vara r�ttsligt bindande .
eldr har f�ljaktligen inte st�llt sig bakom inf�rlivandet av stadgan om de grundl�ggande r�ttigheterna , eftersom r�ttigheterna omfattas av nationell lagstiftning och av europeiska konventionen om m�nskliga r�ttigheter .
men dessa tolkningar , som g�rs av 15 domare och som �verskrider f�rdragen s�som de har ratificerats , �r enligt v�r mening uppenbart lagstridiga . och vi v�ntar fortfarande p� att de skall f� ett godk�nnande fr�n medlemsstaternas folk .
vi borde inte acceptera det , oavsett varifr�n ett s�dant ordval kommer , om det s� �r fr�n extremh�gern eller extremv�nstern !
- ( pt ) de socialistiska ledam�terna fr�n portugal har r�stat f�r duhamels bet�nkande om f�rdragens konstitutionalisering , framf�r allt f�r att de st�mmer �verens med europeiska unionens behov att f�renkla och organisera de grundl�ggande texter som styr den , vilka i dag �r n�st intill ol�sliga med tanke p� den komplexitet som undan f�r undan har ackumulerats i f�rdragen .
den �r i sig �nskv�rd , men antagandet av en s�dan konstitution kan inte vara n�got annat �n en full�ndning av en djupg�ende institutionell reform .
jacques delors har med r�tta p�pekat - f�r knappt en m�nad sedan , bl.a. vid ett sammantr�de i utskottet f�r konstitutionella fr�gor - att termen " konstitution " b�r p� en viktig tvetydighet .
jag skulle till och med r�sta emot , om inte det vore ett alltf�r radikalt s�tt att bed�ma en s� viktig text som denna p� ...
. ( en ) storbritanniens labourledam�ter i pse-gruppen v�lkomnar detta bet�nkande , utan att godk�nna alla dess detaljer .
alla vi vet att europa - dess valuta , diplomati , s�kerhet , civilisation , kultur , sociala modell - inte riktigt kommer att �verleva den lysande historien , men inte heller folkens fruktl�sa kluvenhet , om det inte blir en federation av nationalstater med starka , samst�mmiga och respekterade institutioner som f�reskrivs i en europeisk konstitution , n�got som v�r kollega duhamel m�jligg�r .
avskaffande av villkoren om att ett n�rmare samarbete inte f�r p�verka f�rdragens ramar och avskaffande av vetor�tten och m�jligheten att ta upp fr�gan i europeiska r�det , �r ett brott mot de grundl�ggande principer som det europeiska samarbetet i eu vilar p� .
�ven om bet�nkandet syftar till att i viss m�n luckra upp det mycket rigida system som f�reskrivs under avdelning vii i eu-f�rdraget fr�n amsterdam , vilket �r positivt , �r slutresultatet fortfarande h�gst otillr�ckligt .
europa har faktiskt f�tt det allt sv�rare att g� fram�t med alla medlemsstater .
det �r sk�let till att den omfattande tilldelningen av medel genom eu : s strukturfonder inf�rdes .
om det visar sig n�dv�ndigt med ett f�rst�rkt samarbete �r jag �vertygad om att endast gemenskapssystemet erbjuder de n�dv�ndiga garantierna i form av demokratisk kontroll , r�ttslig kontroll och solidaritet .
vi beklagar ocks� att man inte h�nvisar eller ens n�mner kravet p� att f�rsvara den biologiska m�ngfalden , som �r en av de yttersta randomr�denas viktigaste tillg�ngar .
bryssels europa har - berusad av utj�mning och likriktning - varit or�ttvist och till och med enfaldigt gentemot v�ra medpatrioter , som h�ller v�ra v�rderingar vid liv tusentals kilometer fr�n paris , madrid eller lissabon .
nederl�nderna och danmark har b�da tv� omr�den var i eller p� andra sidan av atlanten men de omr�dena r�knas inte till europeiska unionen .
en av de viktigaste punkterna �r den europeiska livsmedelsmyndigheten . vi gl�der oss s�rskilt �t att den inr�ttas , och vi f�rv�ntar oss mycket av den .
det �r n�dv�ndigt att vi uttrycker oss om ett s� pass viktigt �mne f�r unionsmedborgarna .
detta �r inte alls vitbokens inriktning , eftersom den vill g�ra den europeiska myndigheten till " ett vetenskapligt kunskapscentrum f�r hela unionen " ( sidan 5 ) .
men det �r n�dv�ndigt att g� l�ngre .
f�r min del , i frankrike , har jag inte behov av n�gon myndighet f�r att �terst�lla mitt f�rtroende . jag har f�rtroende f�r afssa ( franska livsmedelsverket ) och dess yttranden , i synnerhet n�r det g�ller galna ko-sjukan .
samtidigt som jag respekterar folks demokratiska r�ttighet att l�gga fram �ndringsf�rslag , m�ste jag �nd� varna kammarens ledam�ter att om vissa av �ndringsf�rslagen som inte finns med i det allm�nna ramavtalet mellan grupperna r�stas fram , s� kommer vi att b�rja �verskrida taken och d�rmed m�ste vi avbryta omr�stningen .
det samma g�ller budgetpost b3-306 f�r informationsprogrammet prince .
det �r ett �ndringsf�rslag fr�n den liberala gruppen om att h�ja tobaksst�det med 5 miljoner euro .
fru talman ! d� m�ste vi tyv�rr r�sta nej till budgetutskottets �ndringsf�rslag s� som det f�rel�g i budgetutskottet .
( parlamentet antog resolutionen . )
bet�nkande ( a5-0270 / 2000 ) av moreira da silva f�r utskottet f�r milj� , folkh�lsa och konsumentfr�gor om kommissionens meddelande till r�det och europaparlamentet om eu : s strategier och �tg�rder f�r att minska utsl�ppen av v�xthusgaserp� v�g mot ett europeiskt klimatf�r�ndringsprogram ( eccp ) ( kom ( 2000 ) 0088c5-0192 / 20002000 / 2103 ( cos ) )
i st�llet f�r att kontrollera de flyktiga kapitalr�relserna prioriteras " strukturreformer " som i sj�lva verket siktar till att privatisera och avreglera sektorer som skulle kunna bli det �nnu mer .
vi menar att medel till balkan i st�llet kan tas fr�n de program i kategori 4 som i dag tyv�rr inte utnyttjas till fullo .
bet�nkande ( a5-0300 / 2000 ) av haug
vi vill ocks� tacka parlamentet f�r den �ppenhet man visade inf�r ett initiativ som enligt v�r mening verkligen f�rtj�nar att uppm�rksammas av denna f�rsamling .
det �r intressant att notera att eu-partierna tydligen inte kan f�rm� vare sig sina medlemspartier eller de enskilda medlemmarna i medlemspartierna att betala en avgift f�r medlemskapet i eu-partiet , utan att man tvingas genomf�ra finansieringen av eu-partierna med offentliga medel .
tilltr�det till accessn�t tvingar n�mligen de offentliga operat�rerna att snarast m�jligt l�mna en prisoffert p� lokalisering av offentliga telefonlinjer .
men : eftersom det handlar om accessn�t m�ste s�rskild h�nsyn tas till kundens intressen .
fr�gan om kvoterna och tr�skelv�rdena kan liknas vid att komma ur askan i elden och det �r en f�r�ndring till det s�mre .
nu n�r det av bilaga iii framg�r att v�xthusodlingen inte drar n�gra f�rdelar av det f�reslagna bidragssystemet f�r gr�nsaker och frukt drar jag tills vidare tillbaka mina inv�ndningar .
" det �r d�rf�r som jag , �ven om jag godk�nner detta dokument , i min r�stf�rklaring understryker att n�sta g�ng skulle det vara l�mpligt att kontrollera och reflektera �ver hur de �ldre och pension�rerna lever i hongkong j�mf�rt med de �ldre och pension�rerna i den folkrepubliken kina , f�r att se om �terf�reningen har varit till gagn eller till skada f�r dem .
bara tre �r har g�tt sedan konferensen i kyoto och europeiska milj�byr�n uppskattar att om utsl�ppen i eu forts�tter i nuvarande takt kommer man inte att uppn� en minskning p� 8 procent av utsl�ppen koldioxid under tiden 1990-2010 utan det kommer i st�llet att bli en �kning p� 6 procent , medan i usa prognoserna �r �nnu s�mre .
f�redraganden anser med r�tta att europeiska kommissionens ursprungliga f�rslag �r otillr�ckligt .
d�rf�r �r v�r resolution som jag har r�stat f�r viktig .
som alla k�nner till �r hela livet genomsyrat av risker och os�kerheter .
vidare b�r en mer konkret ram fastst�llas g�llande forskningen , formaliseringen av tester och samarbetet mellan olika vetenskapliga grupper f�r att uppn� tillf�rlitliga resultat .
vi m�ste g� l�ngre .
de beh�ver i detta sammanhang hj�lp av medlemsstaterna .
h�rigenom skulle dessa f�retag kunna etablera sig fritt inom hela europeiska unionen , �ven om det inte �r n�gra banker .
det �r de �n i dag , f�r alla klagom�l som framf�rs av sm� och medelstora f�retag , missn�jet bland medborgarna �ver h�ga �verf�ringsavgifter f�r mindre betalningar �r fortfarande aktuella .
i praktiken r�cker det med stickprov .
acceptansen av euron �r framf�r allt beroende av om konsumenter och f�retag �r i st�nd att anv�nda euroomr�det som en intern betalningszon .
kanske , nej jag skulle vilja s�ga givetvis , har det blivit tid f�r en internetbank som inte tar ut n�gra kostnader .
fru talman , det finns ett andra sk�l till europaparlamentets ih�rdighet . i bet�nkandet av peijs anges det i sk�l d i resolutionsf�rslaget .
i morse n�dde euron nya bottennoteringar .
i dag uppg�r avgifterna f�r en utlands�verf�ring av 100 euro inom unionen till i genomsnitt 17,10 euro , ett m�ngdubblande av avgifterna f�r inrikes betalningar .
p� sikt f�r det inte finnas n�gon som helst skillnad l�ngre mellan en gr�ns�verskridande och en inrikes betalning .
i denna rapport , s�ger jag nu direkt till peijs i synnerhet , kommer lagstiftningsf�rslag att l�ggas fram om �ndring av det direktiv fr�n 1997 som tr�dde i kraft f�rra �ret .
parlamentet �r i sin vishet helt �verens med er .
sm� och medelstora f�retag �r inte multinationella f�retag i miniatyr , inte heller r�cker det vidare att kvantitativt extrapolera sm� f�retags sv�righeter f�r att uppfatta stora enheters problem p� r�tt s�tt .
fram tills f�r inte s� l�nge sedan f�rest�llde sig de unga att de efter sina studier , efter sin utbildning , antingen skulle s�ka statlig tj�nst eller tj�nst p� ett st�rre statsliknande f�retag .
herr talman , herr kommission�r , k�ra kolleger ! i min egenskap av ledamot sedan elva �r �r jag bland dem som vet att debatter om sm� och medelstora f�retag i parlamentet vare sig �r nya eller s�llsynta .
framf�r allt vill jag i dag pl�dera f�r att l�ta s� m�nga som m�jligt , om inte alla , hinder f�r ett f�rverkligande av den inre marknaden f�rsvinna systematiskt f�r att optimera de sm� och medelstora f�retagens konkurrenskraft , s� att de kan forts�tta att vidareutvecklas p� ett dynamiskt och h�llbart s�tt .
de har den st�rsta anpassningspotentialen .
parallellt f�resl�r vi att ett europeiskt innovationsomr�de uppr�ttas och jag �r f�redraganden tacksam f�r att hon har accepterat att innefatta detta f�rslag i sitt bet�nkande .
vi inst�mmer med den uppm�rksamhet som f�redraganden , montfort , med r�tta �gnar sm� och medelstora f�retag samt mikrof�retag , liksom beviljandet av prioriterat st�d �t unga f�retagare i startskedet .
min partner �r f�r mig specialisten , och n�r jag har n�got problem p� st�domr�det , ett problem med de europeiska institutionerna , kan jag s�ga till mina f�retagare att d�r sitter det n�gon som �r beh�rig och som vet , som p� kort tid kan ge information om offentlig upphandling , om st�dprogram , om forskning kring infrastruktur .
d�rf�r b�r vi vara angel�gna om att med en sn�vare lagstiftning om slim benchmark och best practices s�nka skattesatserna s� mycket som m�jligt f�r att f� enkla och bra regelramar f�r v�ra f�retag .
jag p�minns om vad kommission�ren sade till oss f�r ett �r sedan om sin amerikanska erfarenhet , d�r de inte �r r�dda f�r att misslyckas och tror p� det gamla skotska tales�ttet : " om du inte lyckas direkt , f�rs�k igen och igen " !
i m�nga av v�ra femton medlemsstater har den som �r egenf�retagare j�mf�rt med den privatanst�llde en l�gre niv� p� sin pension , sjukf�rs�kring och f�rs�kring mot arbetsskador .
d�rf�r m�ste vi t�nka " sm�tt " f�rst , " think small first " .
� andra sidan , m�ste vi noga diskutera vilken niv� av europeisk f�rvaltning som �r b�st anpassad f�r det ena eller andra initiativet .
. ( el ) herr talman ! i slutsatserna fr�n europeiska r�dets m�te i tammerfors betonades n�dv�ndigheten av att samarbeta med migranternas och flyktingarnas ursprungs- och transitl�nder och p� uppdrag av r�det utarbetade h�gniv�gruppen f�r asyl- och migrationsfr�gor i samband d�rmed sex handlingsplaner , bl.a. f�r albanien och angr�nsande omr�den .
i mitt bet�nkande har jag tagit alla dessa problem i beaktande och f�resl�r bl.a. : en successiv till�mpning av de �tg�rder som f�resl�s i handlingsplanen , en utredning , som den som g�rs i f�rsta delen , av behoven och som visar p� vilka problem som �r mest akuta , t.ex. m�ste f�rst ekonomin och de demokratiska institutionerna utvecklas , infrastruktur m�ste utvecklas i albanien och d�refter skall unionen forts�tta genom att underteckna avtal om �terv�ndande av flyktingar och migranter .
herr talman ! i handlingsplanens analys fastst�lls att status quo i albanien �r orov�ckande .
( appl�der )
ju t�tare gr�nser vi f�rs�ker skapa , desto vanvettigare flyktingsmuggling kommer vi att f� se .
m�nniskorna hoppas naturligtvis p� en b�ttre politisk representation , men nu finns det fortfarande m�nga m�nniskor som g�r omkring och �ngslar sig , med r�dsla f�r allt och lite till och med r�dsla �ven f�r de v�ldsutbrott som d� och d� f�rekommer .
det finns arbeten t.ex. i grekland som inte skulle kunna utf�ras om de albanska invandrarna f�rsvann , huvudsakligen inom jordbrukssektorn .
det finns f�r n�rvarande en stark str�m av �terv�ndande flyktingar d�r bristen p� s�kerhet , r�ttvisa och ordning st�r i v�gen .
med handlingsplanen som ber�r albanien och angr�nsande omr�den kan man �ka stabiliteten inom omr�det .
p� grund av allt detta , och �ven med anledning av de oacceptabla h�ndelserna i himar , anser jag oss vara tvingade till en mycket f�rsiktig bed�mning av albaniens m�jlighet och vilja att anta de fastst�llda europeiska kriterierna inom omr�dena f�r de m�nskliga r�ttigheterna och de demokratiska friheterna , och f�ljaktligen b�r vi p� motsvarande s�tt �verv�ga och till�mpa v�r allm�nna uppfattning , v�ra handlingsplaner och v�rt bist�nd av olika slag gentemot detta land tills det reviderar sin politik .
en sak till vill jag s�ga .
r�det ( allm�nna fr�gor ) godk�nde redan i oktober f�rra �ret de fem f�rsta handlingsplanerna som g�llde somalia , sri lanka , afghanistan , marocko och irak .
faktum �r att vi har f�rt en mycket seri�s och �ven sj�lvkritisk debatt om kvaliteten p� den europeiska lagstiftningen och till�mpningen av subsidiaritetsprincipen .
vi ber uttryckligen kommissionen ta h�nsyn till den tydliga ansvarsf�rdelningen s�v�l mellan eu och medlemsstaterna som inom institutionerna .
herr talman , herr kommission�r , kolleger ! jag skulle f�rst och fr�mst vilja tacka f�redraganden , wuermeling , f�r det s�tt som han har arbetat med sitt bet�nkande p� .
vi kan acceptera denna �sikt och bet�nkandet �terspeglar andemeningen i detta , genom att man kr�ver en tydligare lagstiftning , en enklare lagstiftning och en proportionerlighet hos de r�ttsliga medlen i f�rh�llande till det efterstr�vade allm�nna m�let .
vi skulle egentligen �nska att kommissionen gav oss fler detaljer om till�mpningen av denna princip med varje f�rslag f�r att g�ra en ordentlig kartl�ggning i samband med �rsrapporten .
maccormick bekr�ftar - och det st�mmer ocks� - att jag sade att subsidiaritetsprincipen inte var en juridisk princip utan en politisk princip .
om staten �r en garant , men ingen h�rskare , s� f�ljer av detta omedelbart att i den konstruktion som gjorts av wuermeling , som i subsidiaritetens namn vill �verl�mna det som i slut�ndan skall garanteras till de enskilda medlemsstaterna , s� m�ste exakt samma process f�ljas �ven av medlemsstaterna .
det �r redan flera talare fr�n europeiska folkpartiets grupp och europademokrater som har framf�rt gruppens �sikter .
det var inte en ordningsfr�ga , utan jag tror att ni i egenskap av f�redragande kunde uttala er f�r att klarg�ra denna fr�ga .
detta direktiv skulle kunna omfatta 64 sidor , vara oerh�rt detaljerat och matematiskt , och involvera m�nga tekniskt sakkunniga .
och
den gamla v�xelkursskillnaden mellan k�p och f�rs�ljning har ersatts av en fast avgift per kontantuttag .
enligt f�redragningslistan f�ljer muntlig fr�ga ( b5-0546 / 00 ) av varela suanzes-carpegna f�r fiskeriutskottet till kommissionen om l�get i f�rhandlingarna om ett nytt fiskeavtal med marocko .
emellertid , n�r detta har sagts , vidh�ller vi ocks� att vi inte godtar vilket avtal som helst .
i v�ra �gon �r det oerh�rt viktigt att gemenskapens fiskare �terupptar sina aktiviteter p� en niv� som �r f�renlig med skyldigheten att s�kerst�lla h�llbara resurser .
som ledamot fr�n den tyska kusten kan jag s�tta mig in i hur fiskarna och deras familjer m�r , som bokstavligen sitter p� torra land , och det sedan m�nader tillbaka .
vi visste alla fr�n f�rsta b�rjan att det var en sv�r f�rhandling .
avtalen med tredje land har en mycket stor betydelse f�r unionen , och i synnerhet f�r regioner med stora fiskehamnar .
det m�ste till grundl�ggande f�r�ndringar , s� att det globala fisket minskar och s� att en mindre del av fiskebudgeten anv�nds till avtal med tredje land .
och jag f�rst�r den europeiska sidan lika v�l : den h�r fr�gan st�r i samband med partnerskapet mellan europa och medelhavsomr�det .
kammaren har varit mycket kritisk mot kommissionen , och det med r�tta , i fr�ga om avtalet med marocko som �nda fr�n b�rjan st�lldes inf�r m�nga oklarheter och naivitet .
herr talman ! herr fischlers fr�nvaro som �r befogad , vilket ordf�randen f�r fiskeriutskottet har understrukit innan , hindrar mig fr�n att g� in p� allt f�r mycket detaljer .
detta inneb�r ett upph�rande av hamnaktiviteterna , fartygsrepareringen , fastygens provianteringsverksamhet , konservfabrikerna , oljefabrikerna , det vill s�ga , att en hel ekonomisk sektor f�r tillf�llet �r lamslagen som konsekvens av detta .
genom detta avtal har n�ra 500 fartyg i europeiska unionen , varav 50 portugisiska fartyg , haft tilltr�de till de marockanska vattnen genom ett �rligt bidrag p� n�ra 125 miljoner euro .
den tillg�ngliga informationen �r knapph�ndig och otydlig , �ven om f�rhandlingarna har fortsatt , s�gs det , med flera besv�rliga f�r�ndringar .
man m�ste skydda v�rldens fiskbest�nd .
men vi m�ste ocks� ha fullst�ndigt klart f�r oss att f�rbindelserna mellan europeiska unionen och de �verg�ngsstater som ligger vid eu : s gr�nser , och till dessa r�knar jag framf�r allt nordafrika , turkiet , ryssland , som �vertar funktionen som �verbryggare mot andra v�rldsdelar och mot andra kulturer vid gr�nserna till europeiska unionen , att dessa stater beh�ver v�rt s�rskilda st�d .
han fick ett positivt intryck av dem , vilket kan ge oss anledning att �nska att de f�rhandlingar som skall inledas den 30 oktober framskrider i en konstruktiv anda .
hj�rtligt tack �nd� f�r detta mycket intressanta bidrag !
texten skulle d� lyda : " att i sk�len ta med att de ber�rda , som �r medborgare i unionen , i hundratals processer i tolv �r varit inblandade i l�ngvariga och upprepade tvister , och att deras ber�ttigade f�rv�ntningar har kommit p� skam .
vi har haft en omfattande skriftv�xling med ber�rda parter och gjort stora insatser f�r att v�lja ut - i h�garna med icke-relevanta dokument - element som p� ett avg�rande s�tt bevisar att de tidigare lettori faktiskt diskriminerades av vissa italienska universitet n�r det g�ller f�rv�rvade ekonomiska r�ttigheter , s�som l�ner och inbetalade avgifter till pensionssystemet .
enligt de italienska reglerna blir man inte universitetsl�rare ope legis , man g�r ett offentligt prov .
om kommissionen vore helt seri�s n�r det g�ller att l�sa denna fr�ga , skulle den ha l�sts f�r flera �r sedan .
det �r inte s� m�nga ledam�ter n�rvarande , eftersom det �r fredag f�rmiddag , men man m�ste notera och inse att detta �r en fr�ga som r�r alla partier och hela unionen .
p� ett kafkaliknande s�tt gick universiteten t.o.m. s� l�ngt att de tog bort l�rarnas namn fr�n de interna telefonlistorna , d�rrarna och universitetens webbplatser .
jag anser att denna mening passar i sammanhanget : " den som inte tar sig sj�lv p� allvar , den blir heller inte tagen p� allvar .
vi inv�ntar en ny dom fr�n europeiska gemenskapernas domstol om den sidan av problemet . det r�r sig s�ledes om tv� saker , som jag inte skulle vilja beskriva som olika , men som �nd� skiljer sig lite �t tidsm�ssigt .
det verkliga problemet �r att vi inte kan godk�nna att en lektor , en person som �r mycket duktig n�r det g�ller engelska spr�ket och som kommer till ett italienskt universitet f�r att f�rklara f�r studenterna vilka som �r de engelska termerna f�r att s�ga hj�rtsjukdom , kirurgiskt ingrepp , leversjukdom osv . , f�r samma r�ttigheter som de personer som undervisar i medicin , samma status .
jag f�rklarar europaparlamentets session avbruten . jag �nskar er en trevlig helg !
vi �r f�renade i chocken och sorgen efter de 150 d�dsoffren och delar de anh�rigas sm�rta .
vad g�ller bet�nkandet av ceyhun f�r utskottet f�r medborgerliga fri- och r�ttigheter samt r�ttsliga och inrikes fr�gor har jag tv� anmodanden : en beg�ran av europeiska socialdemokratiska partiets grupp att �terf�rvisa bet�nkandet till utskottet och en beg�ran av gruppen de gr�na / europeiska fria alliansen att uppskjuta behandlingen av bet�nkandet till ett senare sammantr�de .
( parlamentet godk�nde denna beg�ran . ) tisdag :
fru talman ! min grupp har noggrant lyssnat p� f�rslaget .
b ) sammantr�dena den 29 och 30 november 2000 :
jag hade markerat att jag vill uttala mig innan ni avslutade diskussionen om f�redragningslistan .
detta �r ett mycket allvarligt initiativ som tenderar att �terinf�ra censur i italien , �n s� l�nge bara vad betr�ffar skolb�cker men snart kanske �ven p� andra omr�den .
vi st�der ocks� det bindande i rambeslutet , vilket tvingar medlemsstaterna att anpassa sina lagar till det gemensamma resultatet , samtidigt som l�nderna �r underst�llda den r�ttslig kontroll i eg-domstolen .
parlamentet b�r dessutom vara f�retr�tt i europols styrelse och ha ett ord med i laget vid valet av chef f�r byr�n .
sett ur en mer speciell synvinkel avseende kampen mot penningtv�tt kan vi n�mna r�dets direktiv av den 10 juni 1991 som nyligen �ndrades och f�r vilket v�r kollaga lehne var f�redragande .
jag kan bara s�ga att det som kom fram i slut�ndan visserligen var en riktig uppvisning fr�n r�dets sida , men de �ndringsf�rslag som vi lade fram och som beslutades med mycket stor majoritet h�r i parlamentet antogs inte i det stora hela .
n�r det g�ller dessa fr�gor har v�ra f�redragande behandlat s�v�l det protokoll genom vilket europolkonventionen �ndras som den f�rb�ttrade �msesidiga r�ttsliga hj�lpen .
naturligtvis m�ste bek�mpningen ske p� grundval av enhetliga definitioner om vad brott egentligen �r och vilka metoder som skall anv�ndas f�r att den inte skall kunna undkomma fr�n ett land till ett annat , och d� inte endast av processr�ttsliga sk�l .
jag vill uttala mig om karamanous bet�nkande om europol .
vi har redan alldeles f�r m�nga polisstyrkor och vi kommer att f� �nnu fler n�r v�l utvidgningen �r genomf�rd . v�r f�rm�ga att ta itu med den organiserade brottsligheten kommer att bli mycket s�mre �n vad den borde bara .
vi m�ste se till att de oskyldiga offren - jag antar att vi b�r kalla det den indirekta skadan - i kriget mot brottsligheten inte l�mnas f�r att f�rsm�kta i f�ngelse , isolerade fr�n sina familjer .
i kampen mot penningtv�tten kan vi ifr�gas�tta en fr�ga som , l�ngt ifr�n att vara ett privilegium f�r advokater , �r en grundl�ggande best�ndsdel i r�tten till f�rsvar , som i sin tur �r en grundl�ggande del i v�rt europeiska bygge , kultur och identitet .
vi �r de enda h�r som vill ha �tg�rder som verkligen f�rhindrar penningtv�tt , det vill s�ga ett omedelbart avskaffande av banksekretess , handelssekretess , aff�rssekretess , �ppnande av bokf�ringen i samtliga bank- och industrif�retag samt r�tt f�r f�retagens anst�llda och samtliga konsumenter att offentligg�ra varje kapitalr�relse som g�r emot samh�llets intressen .
enligt fn uppg�r den sammanlagda volymen av det kapital som varje �r tv�ttas till 1 000 miljarder dollar .
n�r det g�ller �tagandena i denna fr�ga avser artikeln antingen de personer som �gnar sig �t en viss verksamhet och d� beh�ver den inte diskutera advokater eller andra yrkesm�ssiga kategorier , eller s� �r det faktum att artikeln tar upp " advokaterna " en situation som i sig sj�lv kan hota den yrkesm�ssiga sekretessen , hur mycket man �n specificerar eller begr�nsar den verksamhet det handlar om .
enligt min tolkning �r " omedelbart " mer kr�vande �n att ge en tidsfrist p� tv� m�nader f�r avvisandet av samarbete .
. ( de ) herr talman , herr kommission�r , k�ra kolleger ! det �r ett frihetens pris att den demokratiska r�ttsstaten ofta ligger efter f�r�varna n�r det g�ller �talen .
h�r har det ansvariga utskottet f�ljt mitt f�rslag , och �ven signalerna fr�n r�det �r gl�djande nog positiva .
det �r inneb�rden i v�ra �ndringsf�rslag .
vi kunde inte f� europol eller interpol att g�ra n�gonting i landet , och det fanns d�lig f�rst�else f�r n�dv�ndigheten av att en person f�r en s� snabb till�ng till domstol som m�jligt .
de straffr�ttsliga systemen h�r ju till en nations mest tydliga kulturella uttryck .
det parlamentet har att ta st�llning till i dag �r ett starkt r�ttsligt samarbete f�r att bek�mpa grov organiserad brottslighet .
. ( fr ) herr talman , jag skulle mycket kortfattat vilja b�rja med att hylla gebhart f�r hennes utm�rkta bet�nkande och s�ga att kommissionen kan ansluta sig till praktiskt taget alla delar som har n�rt dess inneh�ll .
men n�r det g�ller eurojust �r det ett n�tverk f�r samordning av de nationella domarnas och �klagarnas verksamhet i syfte att �ka kapaciteten att k�mpa mot alla former av grov brottslighet p� europeisk niv� .
medan det helt klart �r den nya kommissionen som kommer att avl�gga r�kenskap och m�ste st� till svars f�r denna �rsrapport , handlar det i fair-programmet s� att s�ga om gamla synder ur en f�rg�ngen tid .
min fr�ga om detta till kommissionen pekade p� vissa tillv�gag�ngss�tt , men dessv�rre har hittills inget anv�ndbart resultat utkristalliserat sig .
herr talman ! jag v�lkomnar detta bet�nkande av langenhagen och kan med gl�dje st�dja inneh�llet .
i detta sammanhang vill jag g�rna sl� fast att vi med h�nsyn till den mycket stora sakkunskap som kommissionen har , inte kan acceptera att s� m�nga av de saker som vi har antagit i resolutionerna inte har genomf�rts .
mitt tack g�r s�rskilt till fru langenhagen f�r hennes mycket konstruktiva bet�nkande och till ledam�terna i budgetkontrollutskottet samt fiskeriutskottet , i synnerhet f�redragande busk .
men fr�n och med mitt tilltr�dande tog jag ocks� initiativ till att bilda en informell arbetsgrupp som har unders�kt m�jligheterna att f�renkla och f�rb�ttra f�rfarandena , vilket jag redan har haft tillf�lle att tala om inf�r utskottet f�r industrifr�gor , utrikeshandel , forskning och energi .
ansvaret �r givetvis gemensamt . det �r ocks� revisionsr�ttens sak att uppr�tta dessa dialoger , men jag kan i varje fall f�rs�kra er att det finns en konstruktiv vilja hos revisionsr�tten och kommissionens avdelningar , som ocks� delas av parlamentet , att l�sa dessa problem .
det �r ocks� kommissionens vilja och jag v�gar hoppas att vi kommer att kunna arbeta under b�sta m�jliga f�rh�llanden f�r att genomf�ra detta forskningsprogram , som �r absolut n�dv�ndigt p� europeisk niv� , och m�ste genomf�ras enligt b�sta m�jliga effektivitetsregler men ocks� finanskontrollregler .
herr bethell ! det g�ller inte justeringen av protokollet , men jag kan mycket g�rna tala om f�r er att talmanskonferensen r�stade f�r att f�reningen " basta ya " skall f� �rets sacharovpris .
denna stadga ger ocks� uttryck f�r en gemensam v�rderingsgrund f�r alla kandidatl�nder , f�r alla stater som vill ansluta sig till denna europeiska union , och just n�r det g�ller de sociala r�ttigheterna ger den en klar signal till kandidatl�nderna att de skall uppfylla dessa sociala normer .
. ( fr ) fru talman , mina damer och herrar ordf�rande , mina damer och herrar parlamentsledam�ter ! jag vill f�rst av allt l�ta ordf�randeskapets kondoleanser inst�mma i dem fr�n europaparlamentet , med anledning av katastrofen som �gt rum i n�rheten av salzburg , i �sterrike , och s�ga att vi fullst�ndigt delar anf�rvanternas sorg inf�r denna mycket allvarliga olycka .
ledam�ter i er kammare uttryckte bl.a. vid v�r tidigare debatt �nskem�l om att kunna upprepa denna erfarenhet .
totalt sett skulle jag vilja s�ga att denna text definitivt inneb�r det st�rsta kollektiva framsteget n�r det g�ller att bekr�fta de sociala r�ttigheterna , b�de genom omfattningen av de inskrivna r�ttigheterna , och �ven f�r att dessa r�ttigheter f�r f�rsta g�ngen finns i samma text som de civila och politiska r�ttigheterna , vilket p� ett h�gtidligt s�tt visar att samtliga grundl�ggande r�ttigheter �r odelbara .
jag vill f�r �vrigt ocks� p�peka att ordf�randeskapet , och jag tror �ven �vriga institutioner , �r n�jda med den totala st�ndpunkten fr�n den europeiska fackliga samorganisationen , som betonar den koppling som finns mellan stadgan och den sociala dagordningen , och som sammanfattningsvis anger att slutsatsen av konventet , som antagits av stats- och regeringscheferna , utg�r ett viktigt steg p� " v�gen mot ett socialt och medborgarnas europa " .
d�rf�r var det r�tt och riktigt att europaparlamentet gav utarbetandet av en stadga om de grundl�ggande r�ttigheterna i europeiska unionen en framtr�dande plats och bidrog till den p� ett intensivt och konstruktivt s�tt .
det klarg�rs f�r institutionerna , organen och myndigheterna i europeiska unionen vilka r�ttsliga st�ndpunkter de obetingat m�ste beakta och respektera i sitt agerande f�r m�nniskorna i europa .
v�ra regeringar beh�ver i nice uppn� konkreta resultat att erbjuda medborgarna - de institutionella fr�gorna �r viktiga , men som r�dets ordf�rande och kommission�ren mycket v�l vet �r det sv�rt att s�lja dessa till allm�nheten .
f�r vissa �r det en framg�ng , f�r andra �r det i dag en sviken f�rhoppning .
stadgan kan inte vara en bakgrundsfigur f�r det franska ordf�randeskapet f�r att d�lja en d�ende regeringskonferens .
l�t oss se till att inte samma sak h�nder med f�rdraget om grundl�ggande m�nskliga fri- och r�ttigheter .
vi h�ller p� att programmera ett mord p� kommissionen , ett mord som ocks� �r ett sj�lvmord eftersom kommissionen i f�rra veckan inst�mde i r�dets f�rslag .
fru talman ! f�rst ett hj�rtligt tack till min v�n m�ndez de vigo som ledare f�r delegationen , som har bytt med mig , eftersom jag genast m�ste leda en f�rlikning f�r parlamentet .
hur kan man l�ta bli att erk�nna att bakom konceptet med v�rdighet i det tjugof�rsta �rhundradet �r det samtliga odelbara r�ttigheter som vinner ?
fru talman ! stadgan inneh�ller flera v�lkomna punkter .
det �r tr�kigt att churchills och maxwell fyfes parti har kommit dith�n att de s�ger " nej " , nu n�r vi �ntligen f�rs�ker att se till att unionens institutioner inte blir betraktade som bryssels tyranner , utan som personer som enligt artikel 51 �r bundna till �taganden som skall f�ljas av alla unionens institutioner .
det handlar inte om att g�ra en kolumn med positivt och en med negativt , fru talman .
den andra fascinerande aspekten : vi h�ller i dag p� att diskutera en fr�ga - de m�nskliga och medborgerliga r�ttigheterna - d�r unionen inte har n�gon som helst befogenhet .
p� den punkten �r jag helt och h�llet �verens med honom .
n�gon talare sade att vi m�ste g� ut med information om stadgan , ett arbete som kan inledas i detta parlament .
den �r ocks� modern , som kommissionen p�pekar , eftersom den tar upp fr�gor som handlar om bioetik , genetisk modifiering och informationsskydd , s�v�l som tillg�ng till information .
den som ligger l�ngst efter och som �r s�mst utvecklad har �n en g�ng besegrat den som i samh�llet och i institutionerna k�mpar f�r att de grundl�ggande r�ttigheterna skall g�lla f�r alla och bli ett effektivt och r�ttsligt bindande svar p� nya problem , t.ex. riskerna inom vetenskapen , de nya medborgarnas r�ttigheter , r�tten till en sund milj� etc . vi �r d�rf�r �n en g�ng desillusionerade och missn�jda .
men denna stadga syftar klart och tydligt till att utvidga de europeiska folkens allt n�rmare union .
stadgan �r en balanserad och solid grund f�r utvidgningen .
l�t oss ta v�ra r�ttigheter p� allvar , om vi vill att v�ra regeringar skall respektera dem och om vi vill att v�ra domstolar skall garantera dem .
herr talman ! den stadga som ligger framf�r oss f�r godk�nnande �r ett arbete som vi kan vara stolta �ver .
bara fr�n organisationerna inom europeiska fackliga samorganisationen v�ntas 60 000 m�nniskor .
p� kort sikt �r det mycket viktigare att europeiska unionen binder sig vid europar�dets redan befintliga europeiska konvention om skydd f�r m�nskliga r�ttigheter .
l�t oss g� denna v�g !
jag tycker att man utf�rt ett mycket kvalificerat arbete .
men det finns andra effekter , bl.a. p� v�r egen r�ttsordning .
det mest orov�ckande �r den orwelliknande m�jligheten enligt artikel 52 om upph�vande av de grundl�ggande r�ttigheterna n�r europeiska unionens intressen hotas .
i det h�nseendet vill jag betona att det f�r f�rsta g�ngen i ett dokument fr�n europeiska unionen blir fullst�ndigt tydligt att r�ttigheterna som r�knas upp i stadgan till st�rsta delen beviljas alla m�nniskor , oberoende av nationalitet eller till och med r�tt till uppeh�ll .
kommission�ren har just erinrat om i vilken anda denna stadga utarbetats , som om den skulle bli tvingande en dag .
ocks� h�r �r man ambiti�s med stadgan genom att tillk�nnage r�tten till god administration .
de turkiska medborgarna anser att deras intr�de i unionen inte bara kommer att kr�va en sm�rtfri �versyn av deras institutioner och ett delvis �vergivande av en suver�nitet som de �r mycket f�stade vid , utan �ven en radikal f�r�ndring av deras vanor och mentalitet .
. ( fi ) herr talman , herr minister , kommission�r ! i dag debatterar vi tv� bet�nkanden : morillons �r mer politiskt och mitt mer tekniskt .
i det h�nseendet tvivlar jag inte p� att allas v�r vilja att hj�lpa turkiet att g�ra framsteg p� v�gen mot demokratisering kommer att segra .
ordf�randeskapet anser f�r sin del att detta s�rskilda handlingsprogram f�r l�n fr�n eib mycket snart skall kunna antas av r�det , sannolikt redan vid sammantr�det med ekonomi- och finansministrarna den 27 november .
slutligen m�ste jag s�ga att �ven cypernsamtalet ju har �terupptagits inom fn : s ram .
men jag m�ste ocks� s�ga att jag �r �vertygad om att den turkiska regeringen �r fast besluten att ta itu med de n�dv�ndiga reform�tg�rderna .
jag v�lkomnar ocks� de f�rslag som st�llts i det aktuella bet�nkandet om intensifieringen av det parlamentariska samarbetet och det civila samh�llets starkare roll .
ingenting har gjorts f�r att avskaffa d�dsstraffet . n�stan ingenting har gjorts f�r att p� r�ttslig grund starkare f�rankra minoriteter och m�nskliga r�ttigheter , �ven om vissa fn-konventioner har undertecknats .
herr talman ! europeiska liberala , demokratiska och reformistiska partiets grupp v�lkomnar starkt morillonbet�nkandet , som vi anser har utarbetats p� ett skickligt , uppriktigt och kraftfullt s�tt .
ingen h�r , framf�r allt inte jag , nekar till att det f�rekommit ett folkmord av armenier under den sista epoken av det ottomanska riket .
men d�r handlar det inte bara om att uppfylla k�penhamnskriterierna , utan om demokratiska normer , som �nd� �r absolut n�dv�ndiga .
vi �r helt �verens med denna utsaga , men vi konstaterar att europeiska r�dets beslut i helsingfors att bevilja turkiet status som kandidatland inte f�regicks av en n�dv�ndig allm�n och parlamentarisk debatt , vilket ocks� p�pekas i den n�mnda motiveringen .
man kan inte utnyttja folkens v�rdighet .
r�det kommer att tvingas fr�ga sig huruvida det inte har stj�lpt turkiet snarare �n hj�lpt det genom att ge det kandidatstatus .
( parlamentet antog lagstiftningsresolutionen . )
vi har d�rf�r avst�tt fr�n att r�sta .
i l�nder d�r lagstiftningen �r mer gynnsam f�r arbetarna skulle stadgan d�remot kunna vara g�ngbar mot den .
det eventuella antagandet av stadgan vid det f�rest�ende toppm�tet i nice , antingen genom inf�rlivande i f�rdragen eller helt enkelt som en f�rklaring , inneb�r en negativ utveckling .
artiklar som tr�nger in p� staternas befogenheter .
�ven om l�nderna i europa befinner sig i en alarmerande demografisk situation behandlar stadgan familjeproblemen mycket l�tt .
stadgan kommer att engagera europeiska gemenskapernas domstol i en rad politiska beslut , inom omr�den som �r s� m�ngskiftande som arbetsr�tt , flyktingpolitik , invandring och familjer�tt .
och jag skulle f�rvisso personligen ha f�redragit att dess sociala dimension var mycket mer konsekvent !
. ( fr ) jag bed�mer stadgan om de grundl�ggande r�ttigheterna som ett godtagbart framsteg .
metoden med konsensus som antagits av ledam�terna i konventet har , som vanligt n�r enh�llighet kr�vs , lett till en minimistadga d�r utformningen �r fylld av stora brister och tvetydigheter .
ingen r�tt till arbete , utan " r�tten att arbeta " , ingen r�tt till social trygghet eller till en bostad , utan " r�tten till socialt st�d och st�d till bostad " , ingen r�tt till pension eller en minimiinkomst , inget f�rbud mot upps�gningar , utan ett " skydd mot all omotiverad upps�gning " .
till att b�rja med g�r skillnaderna i �vers�ttning mellan tyskan och franskan att fr�gorna om h�nvisningen till " religi�sa " eller " andliga " v�rderingar kvarst�r fullst�ndigt .
till exempel finns inte r�tten till arbete och r�tten till bostad med .
vi m�ste emellertid best�mt st� emot alla kampanjer f�r en r�ttsligt bindande stadga , som bara skulle skapa r�ttslig os�kerhet .
v�r premi�rminister , ahern , sade nyligen klart och tydligt att europeiska stadgan om de grundl�ggande m�nskliga r�ttigheterna �ven i forts�ttningen b�r vara ett politiskt , inte ett r�ttsligt , dokument .
avslutningsvis har den kohandel som denna typ av process oundvikligen leder till resulterat i att begreppet europ�ernas " religi�sa arv " v�gts mot fr�mjandet av den " fria f�retagsamheten " ...
vidare bygger alla dessa texter p� initiativ fr�n medlemsl�nderna , eftersom de sorterar under antingen den tredje pelaren eller artikel 67 i f�rdraget om europeiska gemenskapen , f�r vilket kommissionen inte har n�got initiativmonopol .
enligt marinhos bet�nkande avser man att utvidga principen med �msesidigt erk�nnande av nationella �tg�rder f�r identifiering , uppt�ckt , frysning eller beslagtagande och konfiskering av brottets instrument och produkter , vilken inr�ttats av den gemensamma st�ndpunkten 98 / 6399 / r�ttsliga och inrikes fr�gor 1998 , till att omfatta beslut som fattas f�re domen , s�rskilt de som skulle g�ra det m�jligt f�r beh�riga myndigheter att snabbt agera f�r att skaffa bevis och beslagta tillg�ngar som enkelt kan �verf�ras .
man accepterade att principen om �msesidigt erk�nnande ocks� skulle till�mpas f�r beslut som fattas under f�rberedande �verl�ggningar , i synnerhet n�r det g�ller dem som skulle g�ra det m�jligt f�r de beh�riga myndigheterna att snabbt s�kra bevis och beslagta tillg�ngar som �r l�tta att flytta .
vi v�lkomnar initiativet fr�n det franska ordf�randeskapet som syftar till att f�rb�ttra samarbetet mellan de nationella myndigheter som �r ansvariga f�r att ta itu med penningtv�tten och fastst�lla enhetliga straffsatser .
. ( en ) samtidigt som jag v�lkomnar ett n�rmare samarbete mellan medlemsstaternas polisstyrkor , b�de mellan dessa och genom europol , delar jag f�redragandens oro �ver bristen p� demokratisk ansvarighet inom europol .
men jag vill rikta uppm�rksamheten p� de m�jliga straffr�ttsliga reformer som kan komma att genomf�ras i olika l�nder - s�som spanien med partido popular vid makten - genom att utnyttja ett visst tillst�nd , f�r dessa reformer �r oroande f�r det fria och demokratiska europa .
bet�nkande ( a5-0310 / 2000 ) av langenhagen
herr talman ! om turkiet vore medlem av eu skulle det vara det folkrikaste medlemslandet n�st efter tyskland .
det h�r �r ett samr�dsf�rfarande , men det rimliga vore f�rst�s att det vore ett medbeslutandef�rfarande eftersom dessa beslut faktiskt kan leda till att budgeten m�ste justeras .
d�rf�r lovordar jag frispr�kigheten som generellt k�nnetecknar morillons bet�nkande , trots att jag anser att en mer direkt formulering p� vissa st�llen skulle ge en mer exakt bild av uppgifterna f�r utv�rdering av turkiets v�g mot anslutning .
med tanke p� detta �r det passande att p� ett f�rd�mande s�tt omn�mna det turkiska flygvapnets bombanfall i kentakor samt att understryka och erinra om den turkiska regeringens skyldighet att villkorsl�st st�dja f�rhandlingarna mellan turkcyprioter och grekcyprioter .
n�stan 40 procent av cypern �r ockuperat av utl�ndsk trupp , av turkiska soldater .
d� m�ste vi konstatera - och det visas ocks� i morillons bet�nkande - att detta inte �r fallet i tillr�cklig utstr�ckning .
vi vill hj�lpa dem p� denna v�g , inte hindra dem , och framf�r allt uppfylla v�ra ekonomiska �taganden .
t�nk s� mycket mer �nskv�rt och godtagbart ett m�l med en l�sare sammanknuten gemenskap av nationsstater skulle vara ; en gemenskap med frihandel och som agerar i samf�rst�nd inom ett begr�nsat antal politikomr�den , och t�nk s� mycket enklare det d� skulle vara att anpassa ett land som turkiet .
vi kan bara inst�mma i denna oro , som kommissionen f�r �vrigt p� ett utm�rkt s�tt gjort sig till tolk f�r i sin senaste �rsrapport .
det nya �r partnerskapet inf�r anslutningen , och i partnerskapet inf�r anslutningen finns det ett mycket viktigt konstaterande . d�r s�gs det n�mligen att kandidatlandet skall behandla alla fr�gor som tas upp i l�gesrapporten .
omr�stningen kommer att �ga rum i morgon kl . 11.30 .
det �r allts� inte f�r att situationen �r sv�r i mellan�stern som konferensen i marseille skall s�nka sina ambitioner .
stora projekt erbjuds �ven samarbetet n�r det g�ller kampen mot all slags illegal handel , migration , och f�rst�rkning av r�ttstaten .
i dag n�r vi st�r inf�r marseille �nskar det franska ordf�randeskapet sj�lvfallet att denna medelhavsprioritering f�r unionen skall bekr�ftas , �ven i ekonomiska termer .
det betyder att det inte bara �r en chans till mer handel och f�r�ndringar , utan ocks� i utomordentligt h�g grad ren s�kerhetspolitik . det m�ste vi tydligt informera v�ra medborgare om , f�r att ocks� f� acceptans f�r det .
det �r visserligen sant att bakslag i den f�rebyggande fredsprocessen har saktat ned framstegen i samband med barcelonaprocessen .
n�r det g�ller de m�nskliga r�ttigheterna , f�resl�r vi ett strukturellt f�rh�llningss�tt d�r man granskar l�ndernas resultat under en viss tidsperiod .
r�det antog i juni 2000 i feira en gemensam medelhavsstrategi och efter att ha f�reslagit och uppn�tt en reformering av medaf�rordningen lade europeiska kommissionen nyligen fram ett dokument om en nyt�ndning f�r barcelonaprocessen .
jag menar till och med att i det f�rflutna har fredsprocessen utgjort ett alibi inte bara f�r europa , utan �ven f�r l�nderna i medelhavspartnerskapet f�r att inte v�ga f�r mycket .
allt detta �r oklart .
dessutom borde dr�mmen om fred p� medelhavets b�da sidor utvidgas och uppfyllas snarast .
braudels " tusen medelhav " , de antika samh�llen som i �ratal betraktat varandra med fientlighet fr�n medelhavets ena strand till den andra har i dag en m�jlighet att inleda en gemensam utveckling , som genom styrkan i dialogen och i den politiska viljan skulle kunna bereda v�gen f�r reella m�jligheter till framsteg och ekonomisk och social utveckling .
genom dess kontinuitet kan den ocks� ge det b�sta m�jliga bidraget , en bieffekt men en viktig s�dan , till �terupptagandet av mellan�sterndialogen .
denna konferens kommer att h�llas inom ramen f�r p�g�ende v�ldsamheter och fredskris , till f�ljd av mellan�sternkonflikten , men det �r ocks� s� att sj�lva dess genomf�rande g�r det m�jligt att h�lla l�gan t�nd f�r europa-medelhavsprocessen och att h�lla den tragiska konflikten utanf�r .
kommissionen och r�det s�ger att de vill det .
f�r det andra anser jag att vi ocks� gl�mmer ett annat viktigt tema , n�mligen milj�n .
nu har en f�rordning lagts fram som i mina �gon g�r det m�jligt f�r europeiska unionen att p� ett effektivt s�tt och i tid hj�lpa l�nderna p� v�stra balkan och tillse att eu-medlen anv�nds p� ett bra s�tt d�r .
det �r anledningen till min uppmaning att inom denna f�rordning finna en god balans mellan synlighet , det vill s�ga stora projekt , � ena sidan och � andra sidan �gna fortsatt uppm�rksamhet �t projekt f�r demokrati , �t projekt som har att g�ra med s�kerhet , projekt som f�r det mesta inte �r s� synliga , men som �r desto mer n�dv�ndiga f�r att garantera stabiliteten p� balkan .
herr talman , herr kommission�r ! jag �r medveten om att balkan inte �r ett omr�de som inger mycket optimism .
vi m�ste genomf�ra ett effektivare och mer samordnat bist�nd och koncentrera alla spridda element .
jag tror att vi alla har klart f�r oss att vi bara med smalare och mer effektiva strukturer verkligen kommer att lyckas att ocks� f�r framtiden stabilisera det goda arbete som kosovobyr�n under de senaste m�naderna har kunnat utf�ra .
jag tror att det �r kontraproduktivt , och jag �r s�ker p� att jacques lang kommer att utnyttja alla sina m�jligheter , och om moscovici skulle vara d�r , skulle han kanske ocks� g�ra det .
enligt min mening g�r huvudpriset denna vecka emellertid till ledarna f�r socialdemokraterna i bosnien och inom parentes till befolkningen i slovakien som inte l�t sig lockas i den folkomr�stningsf�lla som oppositionen hade gillrat f�r regeringen , men det �r ett annat kapitel .
�ret kommer att avslutas med , hoppas vi , konsolideringen av demokratin den 23 december , i samband med riksdagsvalet i serbien .
tilln�rmningen till europeiska unionen �r i r�dets �gon n�ra f�rbunden med utvecklingen av det regionala samarbetet .
det franska ordf�randeskapet hade st�llt upp ambiti�sa m�ls�ttningar f�r v�stra balkan som �r p� v�g att uppn�s : utvecklingen av stabiliserings- och associeringsprocessen , antagandet av cards-programmet , antagandet av asymmetriska handelsf�rm�ner f�r att inte tala om de mest framtr�dande gemenskaps�tg�rderna .
ytterligare m�l f�r toppm�tet i zagreb m�ste omfatta ett tillk�nnagivande av gemenskapens program f�r bist�nd och �teruppbyggnad och demokratisering och stabilisering i v�stra balkanomr�det , ett bekr�ftande av det stegvisa uppr�ttandet av ett frihandelsomr�de mellan europeiska unionen och v�stra balkanomr�det , och ett �tagande av l�nderna i regionen att samarbeta regionalt och uppr�tta ett frihandelssystem dem emellan .
det �r n�dv�ndigt .
sedan flera m�nader har bakers uppdrag tv� m�ls�ttningar . det handlar b�de om att f�rs�ka l�sa de sv�righeter som utg�rs av genomf�randet av planen f�r en l�sning , som b�r leda till att en folkomr�stning om sj�lvstyre f�r folket i v�stsahara genomf�rs och om att f�rs�ka uppn� ett politiskt avtal .
herr talman , herr r�dsordf�rande ! jag tror att eu skulle ha ett mycket st�rre inflytande i maghreb om f�rbindelserna med reformprocessen i marocko vore starkare .
vilka diplomatiska initiativ har r�det f�r avsikt att ta f�r att armenien och azerbajdzjan skall kunna n�rma sig varandra , f�r att den bilaterala konflikten skall kunna l�sas och samarbetet mellan l�nderna fr�mjas ?
. ( fr ) jag f�rst�r de synpunkter som framf�rts av de tv� �rade parlamentsledam�terna . jag har inte mycket att till�gga om unionens �tg�rder s�som de genomf�rts .
herr talman ! jag v�lkomnar r�dets svar p� den ursprungliga fr�gan .
den nya lagstiftning som f�rbereds i turkiet om f�rbud mot straffneds�ttning �r n�dv�ndig , men �nnu viktigare �r att muslimska ledare officiellt tar avst�nd fr�n hedersmord som direkt bryter mot islam .
det spelar ingen st�rre roll om hon syndat frivilligt eller ofrivilligt , dvs. blivit v�ldtagen .
den �sterrikiska regeringen �r den ber�ttigade regeringen i ett av europeiska unionens l�nder . man kan godk�nna dess form eller inte .
jag ville bara s�ga att i den h�r fr�gan f�rel�g ingen diskriminering gentemot det ena eller det andra landet .
n�r ni f�rklarar att h�gerextremistiska partier �r f�rbjudna i �sterrike , s� �r det mycket bra . men man kan ocks� fr�ga sig vad som �r eller inte �r extremh�gern .
n�r det g�ller den politiska l�sningen p� cypern som ni h�nvisar till , herr alavanos , kommer denna fr�ga sj�lvfallet att �ven forts�ttningsvis tas upp med turkiet s�som vi f�rbundit oss att g�ra i helsingfors .
eftersom fr�gest�llaren �r fr�nvarande bortfaller fr�ga nr 11 .
mitt svar var inte s�rskilt pr�glat av optimism eller hopp , utan anger framf�r allt en vilja , den fr�n europeiska unionens franska ordf�randeskap , n�mligen att vi vill kunna sluta ett avtal , ett bra avtal .
delegationen har �ven f�rs�kt att fastst�lla en f�rhandlingskalender .
jag har f�tt ett brev fr�n systern till en annan av mina v�ljare , i vilket hon skriver att hennes bror kvarh�llits i f�ngelse sedan den 28 mars 2000 p.g.a. liknande misstankar .
jag vill , mot bakgrund av det faktum att utvecklingen p� oljemarknaderna kr�ver en mer kraftfull politik av eu p� omr�det f�r energi , fr�ga r�det p� vilket s�tt det tror sig kunna minska den europeiska ekonomins beroende av olja .
. ( fr ) de �tg�rder som den �rade parlamentsledamoten h�nvisar till �terfinns i f�rslaget till budgetlag som undertecknades av president clinton den 28 oktober 2000 .
jag erk�nde att �tg�rder vidtagits av den kubanska regeringen f�r att b�ttre inf�rliva landet ekonomiskt i regionen och jag bekr�ftade p� nytt europas �nskem�l om att vara kubas samarbetspartner i denna process .
f�r det andra h�nvisar r�det som pontius pilatus i sitt svar till nato utan att ta st�llning till turkiets provocerande ifr�gas�ttande av greklands suver�na r�ttigheter , ett ifr�gas�ttande som turkiet den h�r g�ngen passade p� att g�ra med anledning av �vningar med nato .
det �r sant att europeiska unionen ofta anklagas f�r att utlova hj�lp till l�nder som drabbats av olika olyckor eller katastrofer men dr�jer s� l�nge med att ge hj�lpen och att f�rverkliga ekonomiska l�ften att antingen intrycket ges att eu �ngrat sina givna l�ften eller att n�r utbetalningen av pengarna kommer �r det alldeles f�r sent .
f�r det fj�rde , vilket �r mycket viktigt f�r oss : det byggs upp nya gr�nser , men det finns de som alltid l�tt hoppar �ver gr�nserna , n�mligen alla kriminella organisationer med sina brottsliga aktiviteter .
med ett s�dant betraktelses�tt anser jag inte att det tj�nar n�got positivt syfte att �ter ta upp fr�gan ang�ende s�tet f�r europeiska byr�n f�r �teruppbyggnad , en fr�ga som avslutades f�r ungef�r ett �r sedan med packs bet�nkande .
vi m�ste vara medvetna om att v�gen till fred i balkan fortfarande �r l�ng och att det finns potentiella krish�rdar som kan leda till att vi halkar tillbaka ner i det f�rflutna .
jag vill koncentrera mig p� f�rordningarna .
70 procent av de anv�nda medlen hade kontrakterats och 43 procent av de kontrakterade medlen hade betalats .
vi tycker att det �r f�rnuftigare att det n�mns d�r �n att skriva in det i artikeln som handlar om villkor .
spr�kanv�ndningen utg�r ytterligare en k�nslig fr�ga .
detta har utgjort bakgrunden till dessa m�ten .
p� det sociala och kulturella omr�det uppm�rksammade ledarna betydelsen av ett b�ttre samarbete inom utbildningssektorn med s�rskilda initiativ f�r att fr�mja en �msesidig medvetenhet , inklusive en f�rb�ttring av samarbetet mellan universiteten och de elektroniska n�tverken mellan skolor .
om man l�ngsiktigt betraktar den politiska och ekonomiska utvecklingen i v�rlden med sina m�nga poler , �r asiens f�rbindelser med europa och omv�nt av central betydelse .
v�rt problem med asem iii �r inte s� mycket vad som har uppn�tts , f�r det �r naturligtvis positivt med projekt ang�ende penningtv�tt , hiv och aids , livsmedelss�kerhet och liknande .
detta �r sk�let till att europeiska unionen ser till att f� de befogenheter som beh�vs f�r att delta fullt ut .
herr talman ! utan tvekan �r de regionala fiskeorganisationerna i dag den b�sta garanten , om inte den enda , f�r f�rvaltning av v�rldens fiskeresurser och b�r vara det i �nnu h�gre grad i framtiden .
det sker �verfiske , f�rorening av v�ra fiskevatten , klimatet f�r�ndras - det har vi f�rst�tt genom konferensen som p�g�r i haag just nu - och den fysiska f�r�ndringen av milj�n skapar ett �kat tryck p� dessa �ndliga resurser .
fortfarande g�ller den starkares r�tt p� �ppet hav .
l�t mig f�rst och fr�mst ta tillf�llet i akt och v�lkomna bet�nkandet och s�ga att hela fr�gan om f�rvaltning , �vervakning och bevarande av fiskebest�nd utg�r ett st�rre problem .
jag uppmanar kommissionen att ta till sig detta .
i fr�ga om varaktigheten f�r genomf�randet av de regionala fiskeorganisationernas beslut h�ller jag med er om att kommissionens slutresultat kan och m�ste f�rb�ttras .
det �r d�rf�r l�mpligt att t�nka sig nya instrument f�r att vara beredd p� varje allvarlig kris som skulle kunna uppst� , trots en mycket h�g konsumtionsniv� inom unionen och v�l utnyttjade exportm�jligheter .
inr�ttandet av en utj�mningsfond skulle avsev�rt p�skynda koncentrationen i den europeiska slaktgrisproduktionen , eftersom risken med st�rre kapitalinvesteringar skulle �verf�ras till den gemensamma fonden .
den l�ser inte sektorns periodiska instabilitet , den bryter med den gemensamma jordbrukspolitikens solidaritetsprincip och utg�r ett klart fall av �ternationalisering och konkurrenssnedvridning .
om alla gemensamma organisationer av marknaden skulle vara s� anti-cykliskt upplagda som den som garot har f�reslagit , eller om alla organisationer av marknaden skulle komma att verka till f�rdel f�r de mindre f�retagen , vilket ju busk just har anm�rkt p� , d� skulle vi ha en annan struktur p� jordbruksf�retagen i europa .
de senast k�nda fallen av bse kommer att f� en produktionsminskning till f�ljd och st�lla allt som tidigare skett i skuggan .
samtliga medlemsstaters deltagande i detta nya system blir obligatoriskt .
jag �r �vertygad om att man med detta instrument skulle f� st�rre stabilitet p� marknaden och att jordbrukarna i europa skulle f� m�jlighet att beh�rska de cykliskt �terkommande kriserna p� ett b�ttre s�tt .
grisk�ttet har genom tiderna - som keppelhoff-wiechert sagt - drabbats av v�ldigt varierande toppar och dalar n�r det g�ller priset .
jag skulle d� , om vi v�ljer en organisation av marknaden och en f�rst�rkning av politiken p� marknaden , hellre v�lja att g�ra producentgrupperingarna b�ttre rustade s� att de st�r starkare p� marknaden , en marknad d�r de som styr efterfr�gan i allt st�rre utstr�ckning g�r samman och allts� f�r en allt starkare st�llning p� marknaden .
men andra l�nder vill obetingat ha en utj�mningsfond , och jag m�ste helt �ppet s�ga till er : om vi nu skulle f�resl� ett obligatoriskt inf�rande av utj�mningsfonden , skulle f�ljden bli att vi kan gl�mma det hela , eftersom vi aldrig skulle f� majoritet f�r det i r�det .
men rubriken heter h�r : " om f�rslaget till r�dets f�rordning om �ndring av f�rordning ( eeg ) nr 2759 / 75 om den gemensamma organisationen av marknaden f�r grisk�tt " .
de olika kapitlen i �rsrapporten g�ller fyra huvudpunkter .
det fanns ocks� m�nga �verf�ringar av anslag f�r strukturfonderna som avsev�rt �ndrade strukturen av budgeten 1999 . vidare fanns det stora skillnader mellan programbelopp och belopp anslagna i budgetplanen och de flesta av strukturfondernas insatser fick lov att planeras om .
av dessa och andra exempel �r det uppenbart att kommissionen hittills inte bara varit l�ngsam med att vidta korrigerande �tg�rder utan att den i synnerhet har problem med att f� �terbetalning f�r belopp som utbetalats osk�ligt .
men jag blir verkligen f�rv�nad �ver att medlemsstaterna p� tullomr�det till exempel v�grar att �ta sig det finansiella ansvaret n�r deras egen f�rvaltning har gjort fel och tullarna d�rf�r inte kan drivas in , och att de sedan inte tar p� sig det inkomstbortfallet utan alla medlemsstaterna tillsammans m�ste ansvara f�r inkomstbortfallet .
n�r det i slutet av f�rra �ret visade sig att de m�l som fr�n b�rjan efterstr�vades med det humanit�ra st�det inte kan genomf�ras med en l�mplig m�ngd kontroll- och bevaknings�tg�rder , beslutade kommissionen att stoppa aktionen , �ven om det fortfarande fanns medel till f�rfogande .
ni sade , fru schreyer , n�r ni tilltr�dde ert �mbete , att ni skulle f�rs�ka �stadkomma detta .
fru talman ! jag vill b�rja med att tacka revisionsr�tten f�r �rsrapporten .
jag skulle �nska att revisionsr�ttens �rsrapport vore mer konkret .
reformen av kommissionen g�r i h�g grad ut p� att g�ra de enskilda generaldirektoraten ansvariga och jag vill fr�ga revisionsr�tten om den har planer p� att i framtiden omstrukturera �rsrapporten , s� att fler kapitel skapas f�r de enskilda direktoraten .
jag skulle allts� vilja be er svara p� det igen .
jag gl�der mig �ver att kommissionen har vidtagit �tg�rder f�r att f�rb�ttra sin f�rvaltningskontroll �ver gemenskapens finanser och att system inf�rs i medlemsstaterna .
kommissionsreformen garanterar inte att det inte skall f�rekomma n�gra oegentligheter i framtiden .
fru talman ! jag �r ocks� tacksam att r�det har �terkommit f�r jag har n�got att s�ga till dem likas� .
kommer ni , herr karlsson , att f�rbinda er att g�ra detta i framtiden f�r bristen p� tydlig information i rapporten g�r det mycket sv�rt f�r oss att s�tta press p� de r�tta omr�dena , p� de v�rsta lagbrytarna .
f�r att uppn� detta till�nskar jag �ven er , fru talman , stor uth�llighet och jag vill tacka f�r de insatser som ni hittills har gjort .
men ni tar inte med det i rapporten och jag �r tr�tt p� att �r efter �r tvingas h�ra att medlemsstaterna �r ansvariga f�r 80 procent och vi endast f�r 20 procent , samtidigt som det inte anges i rapporten hur det egentligen ligger till !
vi m�ste granska det s�tt som r�tten arbetar p� och hur dess oberoende fr�n institutionerna och programmen den �r avsedd att granska kan f�rst�rkas .
men man m�ste konstatera att vi har att g�ra med ett invecklat system .
i vissa fall handlar det om att ett begr�nsat antal l�nder och ett begr�nsat antal ekonomiska akt�rer som direkt tj�nar p� denna politik .
men jag skulle vilja g�ra det v�ldigt klart att ett f�rfarande av detta slag m�ste utvecklas mycket gradvis s� att vi inte f�r en totalt f�r�ndrad metod f�r att j�mf�ra data f�r d� skulle kvaliteten i detta f�rfarande inte uppfylla kraven i enlighet med f�rdraget .
r�tten �r helt �verens med parlamentet att det inte bara �r en fr�ga om reformering av kommissionen eller om att parlamentet skall reformera sitt s�tt att arbeta med budgetkontroll .
jag t�nkte ocks� p� florida i morse , herr van hulten , och jag �r tacksam f�r att jag inte ansvarade f�r granskningen av valprocessen i just den staten .
jag kan ge ett exempel : n�got jag vet inneb�r sv�righeter f�r r�det , men �r viktigt f�r europaparlamentet och som vi st�der fullt ut �r f�rbudet mot export av produkter som bed�ms vara os�kra till tredje land .
jag �r d�rf�r mycket tacksam till europeiska folkpartiets grupp och europademokrater f�r att det i dag har godk�nt dessa �ndringsf�rslag och �ter l�tit dem bli f�rem�l f�r �verl�ggningar i plenum .
vidare m�ste man naturligtvis fr�ga sig hur pass omfattande de nuvarande standarderna i europa �r och hur pass omfattande de europeiska standarderna skulle vara .
vi befinner oss �n s� l�nge bara i f�rsta behandlingen .
vi m�ste nu titta n�rmare p� kopplingarna mellan produkter och tj�nster .
vi st�der f�r �vrigt kommissionens f�rslag n�r det g�ller ut�kningen av direktivets till�mpningsomr�de till att �ven omfatta tj�nster och migrerade produkter �ven om det p� de omr�dena skulle kunna g�ras mycket mer men det blir vi v�l i alla fall tvungna till i framtiden .
avslutningsvis kan man hoppas att kommissionen kommer att f�rs�ka g�ra den g�llande gemenskapslagstiftningen konsekvent och utveckla den s� att den inte bara blir mer �ppen utan ocks� , eftersom den st�r fast , verkligen kan utnyttjas .
detta �r f�rst�s n�gonting positivt .
direktivets anv�ndningsomr�de m�ste avgr�nsas gentemot de talrika produktbest�mmelserna p� nationell niv� och gemenskapsniv� . d�r regleras �ven de samma s�kerhetsaspekterna .
det har gjorts m�nga anstr�ngningar f�r att definiera hur vertikala best�mmelser , som g�ller vissa produktkategorier , samverkar med detta nya horisontella direktiv och klart tillfredsst�llande resultat har uppn�tts .
den g�ller dock inte n�r specifik sektorslagstiftning som t�cker samma aspekt till�mpas .
jag �r mycket glad �ver att rapporten av fru gonz�lez �lvarez godk�nner huvudprinciperna i kommissionens f�rslag .
denna motivering beh�vs f�r att f�rhindra f�r mycket byr�krati .
i �ndringsf�rslag 19 f�resl�s en harmonisering av medlemsstaternas �vervakningsmetoder p� grundval av riktlinjer utarbetade av kommissionen och den r�dgivande kommitt�n .
i �ndringsf�rslagen 30 , 32 , 42 och huvuddelen av �ndringsf�rslag 33 f�resl�s omformuleringar av direktivets nuvarande text som inte �r f�rem�l f�r revidering .
om kontrollerna bekr�ftar att produkten �r s�ker kommer f�rbudet automatiskt att h�vas .
f�rst kan jag meddela att claudio martelli har �verg�tt fr�n de gruppl�sas grupp till tdi-gruppen , det vill s�ga han har bytt fr�n de gruppl�sas grupp till tdi-gruppen .
( parlamentet antog lagstiftningsresolutionen . )
( parlamentet antog lagstiftningsresolutionen . )
det kan vi tyv�rr inte gl�dja oss �t �nnu .
den f�rsening som har uppst�tt n�r det g�ller att till�mpa avtalen kan bara r�ttf�rdigas till en del .
. - ( en ) jag v�lkomnar detta bet�nkande av averoff om ett f�rslag till att bevilja medel till grekland f�r att minska r�nteb�rdan f�r l�n fr�n eib f�r �teruppbyggnad av regionen attica som blev �delagd vid jordb�vningen i september 1999 .
men alla de p�st�enden som r�r lika m�jligheter f�r kvinnor och m�n f�r en brutal belysning i och med det eu-direktiv som till�ter nattarbete f�r kvinnor .
vi skulle g�rna innan beslutsfattandet om detta femte �tg�rdsprogram ha velat granska det fj�rde .
d� denna icke-statliga organisation spelar en integrerad roll i utformningen och genomf�randet av detta program anser jag att integriteten i denna gemenskapens ramstrategi om j�mst�lldhet mellan k�nen kan ifr�gas�ttas och d�rf�r inte kan st�djas .
. ( en ) medan jag st�der detta bet�nkande om allm�n produkts�kerhet �r det viktigt att vi inte g�r f�r l�ngt .
vi st�der den inriktningen fullt ut , liksom de tv� f�rslag till r�dets f�rordningar som ger den en konkret form , men vi kan inte st�dja europaparlamentets �ndringsf�rslag som syftar till att i grunden �ndra p� balansen i systemet till kommissionens f�rdel .
herr talman ! jag har r�stat f�r bet�nkandet , �ven om inte en tillr�ckligt tydlig �tskillnad g�rs mellan kosovo , serbien och montenegro .
. vi st�der inte nya subventioner till svinuppf�dning och r�star d�rf�r nej till bet�nkandet .
garots bet�nkande syftar till att p� vissa punkter f�rb�ttra kommissionens f�rslag genom att f�rs�ka uppn� en kompromiss med r�det , fr�mst ang�ende medfinansiering av fonden .
. ( nl ) marknaden f�r fl�skk�tt �r cyklisk .
denna f�rsamling talar mycket om r�ttigheter - stadgan antogs i g�r- men n�r det g�ller att till�mpa dessa r�ttigheter , om �n inte i praktiken men �tminstone att betona dem , tar denna f�rsamling skr�mmande stora steg bak�t som verkligen inte �r hedrande .
. det �r utomordentligt att europaparlamentet yttrar sig om turkiets framsteg p� v�gen mot anslutning , s�rskilt vad g�ller respekten f�r de m�nskliga r�ttigheterna .
nu n�r de sista vittnena i exil , de sista som �verlevde blodbadet , sakta d�r ut , blir arbetet och skyldigheten att minnas desto viktigare .
och d� infinner sig kanske �n en g�ng fr�gan om landet verkligen vill bli medlem av europeiska unionen , eller om det inte f�redrar att tillsammans med �vriga l�nder i mellan�stern organisera en integrerad helhet , med mycket n�ra band med europeiska unionen n�r det g�ller handel och ekonomi , s�kerhet och stabilitet samt m�nskliga r�ttigheter och demokratiska spelregler .
de l�nderna h�rde tidigare till det turkiska v�ldet och d�r undertrycktes uppror regelbundet med v�ld .
hela den armeniska befolkning som deporterades till mesopotamiens �knar ; de armenier fr�n �stra anatolien som deporterades p� 24 timmar ; de arbetsf�ra m�n som arkebuserades ; de kvinnor , barn och gamla som f�rf�ljdes och fick g� hundratals kilometer till fots , utan v�rd och mat , som r�nades , v�ldtogs och m�rdades p� v�gen ; de armenier fr�n kilikien och v�stra anatolien som deporterades 1915 ; de 600 framst�ende armenier i konstantinopel som m�rdades ; de mer �n en miljon armenier som avr�ttades p� mindre �n ett �r , dvs. n�stan h�lften av den osmanska armeniska befolkningen - dem f�r vi inte gl�mma .
vi var emot �ndringsf�rslagen om den armeniska massakern av exakt detta sk�l .
totalt sett misskrediteras v�ra intressen ; de f�rsvaras inte med den kraft som �r n�dv�ndig , och kommissionen f�r i f�rsta hand agera som polis gentemot medlemsstaterna , f�r att f� dem att till�mpa de obligatoriska beslut som fattats - ibland mot deras vilja - i den regionala organisationen i fr�ga .
. ( fr ) jag skall inte �terkomma till den utm�rkta argumentation som min v�n gallagher utvecklade ang�ende den text som vi har r�stat om , utan i st�llet utvidga debatten till alla de internationella f�rhandlingar d�r v�ra l�nder f�retr�ds av kommissionen .
ett litet �rende v�xte till slut till ett omfattande arbete genom att farligt och ofarligt avfall samlades i ett direktiv .
lyckligtvis sker det tekniska framsteg . de m�ste s�rskilt anv�ndas f�r h�llbarhetens skull .
vi �r �nd� n�jda med denna tredje behandling , eftersom den st�rker villkoren f�r driftstillst�nd .
det tror jag kommer visa sig vara ett viktigt bidrag till f�rb�ttringen av milj�n .
det �r viktigt att vi inte ers�tter en oh�lsosam och oh�llbar form av avfallshantering med en annan .
jag �r mycket tillfreds �ver denna framg�ng eftersom det inte var l�tt f�r mig som ny medlem att p�verka direktivets andra behandling .
offentlig tillg�ng till information har f�rb�ttrats .
socialf�rs�kringssystemen p�verkas n�mligen av allm�nt utbredda tendenser , som f�r direkta konsekvenser f�r hur de fungerar . det handlar framf�r allt om konsekvenserna av 25 �r med d�mpad tillv�xt , vilket har gett upphov till arbetsl�shet och utslagning samt bromsat skatteint�kterna ; konsekvenserna av befolkningens �ldrande ; konsekvenserna av uppkomsten av nya sjukdomar och slutligen om vetenskapliga och medicinska framsteg som har medf�rt �kade v�rdkostnader .
n�r det g�ller f�ljande punkter skulle det framf�r allt handla om ett f�rslag till rekommendationer : att medlemsstaterna skall erk�nna en gemensam grundl�ggande samh�llsomfattande tj�nst som skall ge alla europeiska medborgare tillg�ng till n�dv�ndig v�rd ; att det i samarbete med de privata f�rs�kringsbolagen uppr�ttas en garanti om att f�lja icke-diskrimineringsprincipen ; att det inr�ttas ett system med �msesidiga f�rs�kringsformer som g�r att kostnaderna f�r omh�ndertagande av personer och grupper med sv�ra sjukdomar delas samt en uppmaning till de privata f�rs�kringsbolagen att utveckla f�rebyggande �tg�rder .
den nuvarande moderniseringen av den sociala tryggheten har som viktigt m�l att garantera ett betalbart h�lsoskydd .
det r�knas som ett socialt europa och det b�r skilja oss fr�n andra .
men varje land f�r sj�lv ta st�llning till vad som �r att f�redra .
jag v�nde mig d� till sjukv�rden och fick beskedet att jag m�ste v�nta tre veckor p� en unders�kning och sedan ytterligare minst en m�nad p� den operation som var alldeles n�dv�ndig .
om alltfler europ�er b�rjar anv�nda till�ggsf�rs�kringar f�r att f� ers�ttning , f�rblir den �msesidiga sektorn den b�sta garantin f�r lika tillg�ng till v�rd .
det g�r nu att �terfinna i fr�mst sk�l j och punkterna 11 e ) och f ) och 14 i det h�r bet�nkandet .
jag tror ocks� att den �kade arbetsr�rligheten i europa beh�vs och ger ett extra argument f�r att l�gga fram en gr�nbok och vidta �tg�rder i fr�ga om sjukv�rdskostnaderna .
men framf�r allt riktar han uppm�rksamheten , till exempel i punkt 3 , p� de betydande problemen med l�ngsiktig h�llbarhet i de allm�nna h�lsov�rdssystemen i hela eu p� grund av de �kande kostnaderna f�r framsteg med behandlingsalternativ liksom det �kande behovet fr�n en allt �ldre befolkning .
mot denna bakgrund anser jag det l�mpligast att vi f�r denna kommissionsunders�kning just om det amerikanska systemet och om systemen i andra l�nder , s� att vi f�r en klar uppfattning om allt detta .
jag m�ste s�ga att �mnet tv�rtom tvingar mig till det , f�r ni , herr talman , framst�r som en �verl�kare med vit rock , stetoskop och hammare att sl� patienterna p� kn�na med .
f�r att undvika missf�rst�nd vill jag �n en g�ng betona att det aktuella bet�nkandet g�ller den kompletterande sjukf�rs�kringen och inte sjukv�rden som s�dan , �ven om det �r s� att de tv� inte f�r skiljas �t .
det �r ett klassiskt exempel p� socialistisk interventionism .
dessa siffror �r dock n�got missvisande eftersom b�de systemens principer och t�ckningsgrad skiljer sig avsev�rt fr�n land till land .
�ven om det r�der stora skillnader mellan de olika medlemsstaterna har portugal den allvarligaste situationen d�r n�ra 24 procent av befolkningen befinner sig i en fattigdomssituation som beror fr�mst p� l�ga l�ner , os�kra och d�ligt betalda anst�llningar och l�ga pensioner som inte ger minsta dr�gliga livsvillkor , varken f�r arbetstagarna och deras familjer , eller f�r �ldre personer .
klagom�l om det fr�n kommissionens sida �r enligt parlamentet ogrundade om det tekniska st�det tas med i sj�lva programmet .
uppdatering av stabilitetsprogrammen f�r tyskland , finland och nederl�nderna
det �r fler och fler medlemsstater som uppn�r en balanserad budgetsituation eller en situation som till och med �r positiv , uttryckt i budgettermer .
i nederl�ndernas fall �r kommissionen bekymrad f�r andra saker , som exempelvis �verensst�mmelsen med policy mix , och de risker som har samband med effekterna av stimulans�tg�rder i form av skattes�nkningar i en konjunktur med en stark ekonomisk tillv�xt , som i nederl�ndernas fall skulle kunna ge upphov till en �verhettning .
herr talman , herr kommission�r ! herr kommission�r , vi �r tacksamma f�r den rapport ni har avlagt om utvecklingen av den nya nettoskulden i europeiska unionen .
herr talman ! jag tycker ocks� att det �r h�rligt att se att det sker en positiv utveckling inom de offentliga finanserna i de ber�rda l�nderna , men jag har lagt m�rke till att m�nga m�nniskor i dag �r oroliga f�r hur det skall g� med prisstabiliteten i europa .
jag skulle vilja veta om kommissionen kan ge n�gra upplysningar om detta , herr kommission�r .
europeiska unionens r�d agerar s�ledes aktivt , tillsammans med er institution och europeiska kommissionen , f�r att modernisera och st�ndigt f�rst�rka det europeiska systemet f�r att f�rebygga och motverka denna sjukdom .
kontrollresurserna i hela livsmedelskedjan kommer att f�rst�rkas .
den europeiska livsmedelsmyndigheten skall ocks� tillhandah�lla tydlig och l�ttillg�nglig information i fr�gor som sorterar under dess mandat .
om dessa kontroller beaktas och genomf�rs minskar risken f�r allm�nheten till ett minimum .
kommissionens �sikt att riktad provtagning �r avg�rande f�r att f� en sann bild av den verkliga f�rekomsten av bse i gemenskapen har visat sig vara helt riktig genom provresultaten i frankrike .
specificerat riskmaterial m�ste tas bort och f�rst�ras .
l�t mig till�gga n�gra synpunkter p� det som jag sade tidigare i detta h�nseende .
jag v�lkomnar ocks� i detta avseende att premi�rminister jospin i g�r ocks� meddelade en v�sentlig f�rst�rkning av kontroller i livsmedelskedjan , inklusive en stor personal�kning .
men till�mpningen i medlemsstaterna sker fortfarande alldeles f�r l�ngsamt .
jag vill tydligt p�peka , kolleger , att det vi beh�ver �r tv� saker .
i en situation som den som nu har uppkommit i frankrike , och �ven tidigare i m�nga andra l�nder , �r det angel�get att kunna tala om f�r konsumenterna var de produkter som de f�r kommer ifr�n och hur dessa produkter kan sp�ras .
de som i dag h�vdar att de inte har n�gra fall av bse p� deras territorium , herr b�ge , �r de som inte s�ker efter s�dana fall .
det �r d�rf�r br�dskande att vidta �tg�rder f�r att lugna konsumenterna och �tervinna deras f�rtroende f�r livsmedelsprodukters s�kerhet .
jag skall inte i detalj r�kna upp alla de ohyggligheter som har beg�tts av �n den ene �n den andre .
den franska regeringens �tg�rder �r i det avseendet otillr�ckliga .
en sak som k�nnetecknar d�liga avtal �r att de m�ste ifr�gas�ttas , och sk�len blir s� mycket starkare n�r folkh�lsan kr�ver det .
men i den h�r krisen m�ste vi garantera att s�v�l konsumenternas h�lsa och livsmedel som uppf�darnas inkomster skyddas , det g�ller t.ex. slaktare , f�rs�ljare av in�lvsmat , grossister - alla som fallit offer f�r statsmakternas slarv , s�v�l nationernas som gemenskapens .
fru talman , herr r�dsordf�rande , herr kommission�r ! den h�r debatten har �tminstone f�rdelen att den avsl�jar meningsskiljaktigheterna mellan oss alla , mellan r�det � ena sidan och kommissionen � andra sidan .
en reform av den gemensamma jordbrukspolitiken �r inte bara n�dv�ndig : den �r ofr�nkomlig , eftersom det inte �r godtagbart att endast ett land vidtar str�nga �tg�rder och f�rs�tter sin ekonomi i sv�righeter .
d� skulle man inte nu beh�va klaga �ver att man placeras i en kategori som man inte ville placeras i , eftersom man endast postulerat att ingen bse f�rekommer .
f�r att kostnaderna f�r krisen inte helt skall drabba uppf�darna kr�ver vi att de f�r ekonomisk hj�lp .
jag vill dock p�peka att ingen m�nniska klarar sig utan mat , inte ens en dag .
herr byrne sade inte s� mycket i dag , fast�n han var mycket efters�kt f�r att g�ra det om tester .
f�r det f�rsta : f�r att bem�ta den europeiske konsumentens ber�ttigade och mycket kr�vande behov av livsmedelss�kerhet , l�gger vi ribban mycket h�gt n�r det g�ller kontroller och f�rsiktighets�tg�rder .
till�mpa i st�llet det vi har beslutat , s� beh�ver vi inte diskutera den h�r fr�gan mer .
d�rf�r m�ste konsumenter och producenter f�rena sig f�r st�rre s�kerhet med utg�ngspunkt i den okr�nkbara principen att mat skall vara h�lsosam .
och om vi hade den politiska viljan , kan jag f�rs�kra er att det h�r problemet inte skulle finnas i dag , f�r alla fakta om problemet �r k�nda .
f�r det andra handlar det om att anv�nda benmj�l i djurfoder eller inte , vilket det �ven h�r f�rs en livlig debatt om .
vi ser allt oftare �ven i v�rt land att ett d�tt f�r eller en d�d kalv helt enkelt l�mnas kvar , eftersom det �r f�r dyrt att l�ta h�mta det .
det brittiska systemet att ta bort smittade djur fr�n bes�ttningarna och betala bra ers�ttning f�r dessa djur uppmuntrar b�nder att tillk�nnage sina fall av bse .
kommission�r byrne var mycket kraftfull i sitt �ppningsanf�rande n�r han sade till kammaren att han vara beredd att titta n�rmare p� denna fr�ga om k�tt- och benmj�l och g� vidare med den .
de hj�lper oss att g�ra framsteg , och d�rf�r har jag med stor uppm�rksamhet lyssnat till alla era anf�randen , f�r i det h�r skedet tycker jag att det �r l�mpligt att debatten om unionsmedborgarnas s�kerhet f�rs p� europeisk niv� .
det som vi m�ste komma ih�g n�r vi �verv�ger denna fr�ga �r det faktum att det redan finns ett f�rbud mot att utfodra boskap med k�tt- och benmj�l .
de tester som jag h�nvisar till nu �r n�got olika .
p� grund av den senaste tidens frekventa h�ndelser i olika medlemsstater , d�r de mest grundl�ggande m�nskliga r�ttigheterna inte har respekterats vid avvisningen eller utvisningen av invandrare , b�r denna fr�ga specialgranskas av kommissionen .
herr talman ! jag vill s�ga att jag ansluter mig till fru ledamotens oro och hoppas att era krav inte bara riktas till kommissionen , utan ocks� till r�det , s� att hela den r�ttsliga ramen kan godk�nnas till juni n�sta �r .
vilka �tg�rder �mnar kommissionen vidta f�r att f� ett slut p� denna situation av grovt utnyttjande , misshandel och handel med vita m�nniskokroppar , en situation som absolut inte kan tolereras - och vad �mnar kommissionen g�ra f�r att avskaffa alla former av kvinnodiskriminering ?
kommer kommissionen att vidta n�gon �tg�rd f�r att �tminstone s�tta stopp f�r de m�nga olika �sikter som f�r n�rvarande r�der och som s� allvarligt skadar eurons utveckling ?
jag ber er , ledam�ter , att b�rja med fr�gan och inte med f�rklaringen .
kommissionen har d�rf�r nyligen �verl�mnat ett yttrande till de grekiska myndigheterna .
. ( en ) om v�rdena �verskrids m�ste medlemsstaten , i detta fallet grekland , vidta �tg�rder .
. ( fr ) n�r kommissionen beslutade att godk�nna det franska systemet f�r st�d till filmproduktion , fastst�llde vi fyra specifika kriterier f�r f�renlighet .
vi f�r dock inte n�ja oss med det vi hittills har uppn�tt .
f�r det f�rsta genom att f�rb�ttra f�rst�elsen f�r utslagningen som fenomen , med hj�lp av indikatorer och utv�rderingskriterier , som framf�r allt �r inriktade p� m�lgrupper .
man s�ger till oss att det b�sta s�ttet att f�rhindra social utslagning �r att hitta ett betalt arbete men jag skulle vilja h�lla med dem som har sagt att vi m�ste ta h�nsyn till det faktum att inkomstbringande syssels�ttning inte enbart �r en garanti f�r socialt deltagande .
det kan g�lla �ldre m�nniskor , vars kunskaper inte l�ngre beh�vs .
p� de h�ll i europa d�r detta har gjorts har man uppn�tt best�ende minskningar av arbetsl�sheten .
dessutom lever enligt eu : s statistiktj�nst 18 procent av de europeiska medborgarna under fattigdomsgr�nsen , medan en tredjedel av de som �r fattiga arbetar .
en g�ng om �ret �ker jag tillsammans med mina v�nner thomas mann och mario mantovani till poverelle-instituet i bryssel ; d�r serverar vi mat till de stackars luffarna och v�ra hj�rtan bl�der och vi k�nner skuld �ver att vi bara g�r det en g�ng om �ret . vi skulle vilja g�ra det varje dag , men det kan vi uppriktigt sagt inte .
det �r ett ambiti�st program f�r gemenskaps�tg�rder , enligt kommissionens f�rslag , det kommer att f� 70 miljoner euro i budgetanslag och g�lla under en period p� fem �r .
avslutningsvis vill jag g�rna �terigen sl� fast att solidariteten mellan staterna m�ste vara den grund p� vilken man skall bygga en solid ny kamp mot fattigdom och social utslagning . emellertid m�ste man ta h�nsyn till att de ekonomiska framstegen i medlemsstaterna , och d�rmed deras �kade v�lst�nd , med till�mpning av skalf�rdelarna i den sociala marknadsekonomin s�kerligen kommer att medf�ra att man kan skapa en st�rre och b�ttre social r�ttvisa .
jag h�ller ocks� med om att det �r viktigt att �ka f�rst�elsen f�r social utslagning och fattigdom och att ta fram j�mf�rbara indikatorer och bed�mningskriterier .
men jag skulle vilja ge f�ljande pragmatiska f�rslag som svar p� era farh�gor , f�r jag h�ller helt med om att vi m�ste hitta en metod f�r n�ra och kontinuerligt samarbete .
fr�mjande av el fr�n f�rnybara energik�llor
s� mycket tid har vi inte !
f�r att f�rtydliga det hela : f�rbr�nningen av avfall �r ingen f�rnybar energik�lla och kan d�rf�r inte heller bidra till uppfyllandet av m�len .
vi anser att dessa riktlinjer , om de inte �ndras , kommer att ge upphov till mycket negativa milj�effekter .
kolleger , detta direktiv l�ter vettigt .
efter generaladvokatens pl�dering i eg-domstolen i luxemburg �r risken inte lika stor f�r att prisst�den upph�vs av best�mmelserna f�r statligt st�d .
vi f�rs�ker inte f� andra att tro att torveldning skulle minska koldioxidutsl�ppen , men torven �r ett inhemskt br�nsle , medan olja och gas �r importvaror .
oljan kan inte ers�ttas med kol , naturgas eller uran .
vi �r f�r en kortare period och d�refter en utv�rdering och jag vill s�ga till min kollega , fru mcnally , att hon m�lar en vacker bild av vindkraftanl�ggningar i havet , men jag m�ste s�ga till henne att de tekniska problem och de kostnader som det handlar om g�r att den tekniken , liksom elektricitet fr�n solen , har ganska l�ng v�g kvar tills den kan anv�ndas i framtiden .
naturligtvis pekar detta direktiv i r�tt riktning : n�mligen , �ntligen , ett seri�st v�rdes�ttande av de f�rnybara energik�llorna .
herr talman ! jag vill tacka min kollega roth f�r det v�rdefulla arbete han utf�rde vid utformandet av bet�nkandet .
v�r m�ls�ttning med avseende p� h�llbar energi �r ambiti�s men i samband med klimatproblemen �r vi �nd� blygsamma .
herr talman ! det f�r inte finnas n�gra tvivel om att en kombination av investeringar i f�rnybara energik�llor och energieffektivitet �r det enda realistiska s�ttet f�r europeiska unionen att klara av kraven i kyotoprotokollet och minska v�rt tunga beroende av fossila br�nslen .
vi m�ste med mycket bred majoritet r�sta f�r f�rslagen fr�n rothe .
n�r det g�ller v�ra m�l p� omr�det , m�ste vi lyssna p� medborgarna och str�cka oss l�ngre �n kommissionens f�rslag , som jag betraktar som mycket positivt i sin helhet , p� 21 procent , och �ka den f�rnybara delen av den totala elproduktionen .
i �ndringsf�rslag 1 , 2 , 8 , 20 och 21 understryks behovet av en politik som fr�mjar den gr�na elen och alla f�rdelar med denna och dessa godtas utan vidare av kommissionen .
d�rf�r st�der vi �ndringsf�rslag 36 och 56 och �ven vissa aspekter i �ndringsf�rslag 4 , 15 och 62 , som har att g�ra med tanken p� en internalisering av de externa kostnaderna och kompensationen f�r de uteblivna externa kostnaderna till f�rm�n f�r de f�rnybara energik�llorna .
kvinnors deltagande i fredlig l�sning av konflikter
kvinnor m�ste delta fullt ut i alla fredsf�rhandlingar , i allt �teruppbyggnadsarbete och i fredsbevarande operationer .
kvinnornas situation framst�r dock som s�rskilt sv�r n�r de precis som tidigare m�ste k�mpa f�r ett erk�nnande och ett deltagande p� lika villkor .
det motst�nd som vissa m�n i den h�r kammaren visat mot en seri�s behandling av det h�r �mnet �r ett tydligt tecken .
man kan �ven undervisa om anlitandet av frivilligorganisationer , uppbyggande anordningar f�r krisdrabbade personer etcetera . vi kunde sedan anordna utfr�gningar , seminarier och s� vidare i dessa fr�gor .
vi h�ller med om erk�nnandet att v�ldt�kter , p�tvingade graviditeter , p�tvingad sterilisering och alla andra former av sexuellt v�ld utg�r brott mot m�nskligheten , och d�rf�r b�r lagtexten aktualiseras f�r att ge ett effektivt skydd �t kvinnor .
( talmannen avbr�t talaren . )
mina gratulationer en g�ng till och l�t oss hoppas att det leder till resultat .
i bet�nkandet tas inte bara kvinnors sociala utslagning upp som ett problem i sig utan det po�ngteras ocks� helt riktigt att skyddet mot brottslighet och den personliga s�kerheten inte l�ngre bara kan garanteras inom nationens gr�nser .
p� det h�r omr�det finns det inget annat �n pinsamma misslyckanden och trots detta m�ter vi fortfarande en mur som utest�nger kvinnorna .
i iver att vara emot allt ont f�rd�ms systematiska v�ldt�kter och sexuellt slaveri .
det fj�rde exemplet �r kvinnornas viktiga roll i den av europeiska gemenskapen st�dda fredsprocessen p� balkan och i medelhavsomr�det .
. ( nl ) herr talman ! vi �verg�r nu till ett mer jordn�ra problem , n�mligen enhetliga best�mmelser f�r hush�llsarbete som utf�rs av utomst�ende personer i privata hush�ll , det �r ju det som det handlar om .
slutligen m�ste allt detta n�dv�ndigtvis inneh�lla ett ekonomiskt ingripande fr�n myndigheterna , fiskalt eller parafiskalt , ett privathush�ll kan n�mligen inte betala en fullst�ndig stadga , �ven om den �r begr�nsad , och d� stannar alla kvar p� den svarta marknaden .
arbetstagarna , som huvudsakligen �r kvinnor , b�r f� �kad tillg�ng till utbildning .
herr talman , herr kommission�r !
herr talman , fru kommission�r ! hemhj�lp , n�got som tidigare n�stan enbart anlitades av v�lbest�llda hem , har i dag blivit en n�dv�ndig och oumb�rlig hj�lp f�r yrkesverksamma kvinnor och m�n , och i synnerhet �ven f�r ensamst�ende m�drar och �ldre .
omr�stningen kommer att �ga rum i morgon kl . 12.00 .
vi f�rv�ntar oss mycket av ert anf�rande , herr president ; att ni visar v�gar f�r detta �terfunna samarbete och broderskap , v�gar som vi numera kommer att g� tillsammans . det �r en gl�dje f�r mig att nu ge er ordet .
vi skall inte bara genomf�ra privatisering av v�r centraliserade ekonomi utan ocks� skapa ett r�ttsligt system som skall garantera frihet f�r aff�rsverksamhet och f�r hela den ekonomiska processen .
n�r det g�ller f�rbindelserna mellan serbien och montenegro inom den federala staten hotade den forna icke demokratiska organisationen i den federala republiken jugoslavien allvarligt statens funktion .
d� inledde era modiga f�reg�ngare ett os�kert projekt som gav historiskt resultat .
justering av protokollet fr�n f�reg�ende sammantr�de
herr talman ! mitt �rende g�ller mera framtiden �n det f�rflutna , jag vill n�mligen f�rs�kra mig om att omr�stningen i fr�gan om bse sker i dag .
i b�rjan av denna valperiod l�mnade jag sj�lv in ett fullst�ndigt initiativf�rslag till utskottet f�r konstitutionella fr�gor .
den h�r r�tten b�r naturligtvis avgr�nsas , och �ven detta b�r vi diskutera i dag .
herr talman ! parlamentsledam�ternas r�tt till tillg�ng till sekretessbelagda dokument �r mycket viktig , men den kan inte ers�tta medborgarnas r�tt att f� direkt information .
det �r dessa �verv�ganden som har f�rm�tt budgetkontrollutskottet att avge ett yttrande i detta �rende .
deras kunskaper �r beroende av �sikterna i media eller s�rskilda intressegrupper och de k�nner ofta vanmakt gentemot institutionerna .
nu g�ller fr�gan dock allm�nhetens , inte parlamentets , tillg�ng till handlingar .
vi har d�rf�r minskat dem till 6 .
dessutom skall det varje �r l�mnas en rapport till parlamentet , s� att vi fortl�pande kan f�lja upp denna verksamhet .
begr�nsningarna av kommissionens och r�dets informationsplikt gentemot europaparlamentet h�r inte hemma i detta lagf�rslag .
med andra ord uppr�ttas en , i mina �gon , felaktig l�nk mellan parlamentsledam�ters r�ttigheter och allm�nhetens r�ttigheter .
s� till de punkter d�r vi k�nner os�kerhet : den f�rsta g�ller sektorerna gemensam utrikes- och s�kerhetspolitik , men �ven r�ttsliga fr�gor och inre angel�genheter .
f�rordningen kan principiellt betraktas som positiv , framf�r allt klarg�randet att denna f�rordning omfattar b�de alla politikomr�den och alla institutioner inom unionen .
herr talman och k�ra kolleger ! jag riktar en uppmaning till er om att vi skall f�rs�ka f�rm� r�det att �ndra �sikt och samtidigt riktar jag en uppmaning till er att r�sta f�r cashmans bet�nkande .
herr talman ! jag vill tacka f�redraganden och alla andra som har varit inblandade i detta arbete .
till sist : det existerande hemligh�llandet �r till och med f�r parlamentsledam�terna s� stort att m�nga sammanhang som vi beh�ver k�nna till f�r det egna beslutsfattandet f�rblir s� dolda , att man ...
vi ledam�ter b�r ha mer mod .
det vore b�ttre att skriva in regler som f�rpliktar alla enheter att offentligg�ra och registrera sina handlingar .
denna klyfta symboliserar avst�ndet mellan europeiska unionen och dess medborgare .
jag vill till�gga hur mycket jag och kommissionen uppskattar cashmans och f�rfattarinnan till f�rslaget maij-weggens anstr�ngningar f�r att p� s� kort tid l�gga fram detta bet�nkande .
jag tror att det visar att det inte finns perfekta situationer , och att vi m�ste g� vidare tillsammans f�r att undvika situationer som denna .
h�ri innefattas �ndringsf�rslag som de som presenterats om �tg�rder som man b�r komma �verens om genom interinstitutionella avtal : nr 34 , 45 och 48 .
jag framf�r den h�r synpunkten med tanke p� att den kommission�r som kommer hit vanligtvis ger en muntlig presentation av kommissionens rekommendationer till omr�stning .
omr�stningen kommer att �ga rum kl . 12.00 .
v�rt utskott accepterar kommissionens f�rslag om en extern ratingfunktion , med reservationen att detta �r en funktion med begr�nsningar och att det viktigaste �r att sm�f�retagen inte skall beh�va bli taxerade och inte heller skall f�retag utan taxering bli eftersatta .
( parlamentet antog resolutionen )
bet�nkande ( a5-0318 / 2000 ) av cashman f�r utskottet f�r medborgerliga fri- och r�ttigheter samt r�ttsliga och inrikes fr�gor om f�rslaget till europaparlamentets och r�dets f�rordning om allm�nhetens tillg�ng till europaparlamentets , r�dets och kommissionens handlingar ( kom ( 2000 ) 30 - c5-0057 / 2000 - 2000 / 0032 ( cod ) )
majoriteten av kvinnorna skall resa till en konferens med parlamentariker i berlin .
bet�nkandet av villiers f�rtj�nar b�ttre �n att g� till omr�stning i morgon f�rmiddag .
jag g�r med p� detta , men om ni hade f�ljt f�redragningslistan , och inte f�rst hade l�tit bet�nkandet fr�n cashman g� till omr�stning d�rf�r att ett antal personer inte kommer att vara n�rvarande i kv�ll , f�r detta �r orsaken , s� hade vi �ven kunnat r�sta om smetbet�nkandet .
n�r det g�ller ert f�rsta p�pekande , ledamot mann , s� kommer det naturligtvis att skickas till parlamentets presidium och till talmanskonferensen .
. kommissionen och europeiska unionens r�d har ett stort ansvar f�r den omfattning som fr�gan om bse hos n�tkreatur har f�tt .
vad g�ller inneh�llet har min grupp rekommenderat str�ngare �tg�rder f�r att bek�mpa epidemin .
den tvetydiga formuleringen i punkt 4 kan dessutom bara v�cka fr�getecken kring myndigheternas vilja att med alla tillg�ngliga medel mots�tta sig de agrara livsmedelstrusternas svindel och bedr�gerier , n�r det vore s� mycket enklare att med en enda mening sl� fast att produktion och anv�ndning av animaliskt mj�l �r helt f�rbjudet .
folkh�lsan m�ste vara den gemensamma jordbrukspolitikens fr�msta m�l .
de fall av bse som f�rekommit i frankrike , liksom fallen av dioxinsmittade kycklingar i belgien , �r de senaste i en l�ng rad av f�rsummelser .
wto-f�rhandlingarna m�ste �terupptas , s� att de europeiska jordbrukarna kan �ka sin produktion av proteiner av vegetabiliskt ursprung .
kommissionen planerar synbarligen ingenting annat �n genomsnittliga �tg�rder , vilket inneb�r att de stater som �r mest kr�vande i fr�ga om s�kerhet inte kommer att f� ett " plus " , utan ett " minus " , n�got som i subsidiaritetsprincipens namn b�r vara en anledning till att �terge medlemsstaterna friheten att vidta de �tg�rder som kr�vs f�r att effektivt skydda sina befolkningar och garantera deras s�kerhet , mot bakgrund av opinionsl�ge , politisk vilja , epidemitillst�nd samt den st�llning som de ber�rda sektorerna har i l�ndernas ekonomi och samh�lle .
dessa legitima farh�gor ledde till att parlamentet visade stor uppm�rksamhet och l�mnade in �ndringsf�rslag i syfte att strikt reglera allt som r�r f�rbr�nnings- och samf�rbr�nningsprocessen .
alla dessa �tg�rder avspeglar allm�nhetens f�r�ndrade �sikter om �mnet avfallshantering .
att samh�llsinstanserna och s�rskilt f�retr�dare f�r de utsatta grupperna till vilka programmet �r riktat medverkar i processen ,
det �r min plikt att v�lkomna det h�r initiativet , som bem�ter medborgarnas f�rv�ntningar .
detta kommer att uppn�s genom att st�lla upp specifika m�l som skall integreras i de nationella handlingsplanerna och att genomf�ra en politik f�r att fr�mja lika m�jligheter .
samtidigt som den ekonomiska tillv�xten �r stark och arbetsl�sheten tenderar att g� tillbaka , �r ett arbete i dag inget skydd mot utslagning .
den brittiska labourregeringen har lett kampen mot fattigdom och social utslagning .
det l�mnas miljardsubventioner till n�gra f� som f�rst�r landskapet med sina vindkraftverk .
medlemsstaterna m�ste nu sl� in p� den h�r v�gen f�r att respektera de milj�m�l som de har skrivit under p� , b�de p� europeisk och internationell niv� , men ocks� f�r att s�kerst�lla sitt energioberoende och en s�ker elf�rs�rjning .
d�rf�r �kar k�rnkraftens betydelse hela tiden .
k�rnenergi kan leda till katastrofer som g�r stora delar av v�rlden obeboelig , och producerar en farlig avfallsprodukt .
det �r br�dskande att �teruppliva den interparlamentariska dialogen mellan v�steuropa och �stra asien .
vi anser att den regionala integrationen �r ett avg�rande instrument f�r att fr�mja de tre grundl�ggande m�l som jag har n�mnt .
jag tror att det var fyra �r sedan som vi p� kallelse av irela tr�ffades i antigua , en oerh�rt vacker stad i guatemala . d�r diskuterade vi med v�ra kolleger i det centralamerikanska parlamentet vad det skulle bli i framtiden , inte bara f�r det centralamerikanska parlamentet utan ocks� f�r europaparlamentet .
d�rf�r b�r man enligt mitt s�tt att se det helt och h�llet avvisa den kritik fr�n intresserade parter som beskyller det centralamerikanska parlamentets verksamhet f�r att vara ett konstgjort system eller parlamentarism av tom , ih�lig och inneh�llsl�s papjemach� .
i detta sammanhang agerar kommissionen och p� de tre niv�erna har vi olika projekt .
( b5-0849 / 2000 ) av rod och maes f�r verts / ale-gruppen ;
det �r hela inneb�rden av v�r resolution .
en l�ngvarig fred �r dessutom ot�nkbar i detta land utan religi�s och etnisk tolerans .
men enligt min mening , herr talman , m�ste vi framf�r allt vara mycket beslutsamma n�r det g�ller kravet p� att den rasistiska konstitutionen ogiltigf�rklaras .
�ven han har ju dragit det nationalistiska kortet .
vi kan bara se till att detta blir ett fritt och fredligt val , och hoppas att elfenbenskustens ny regering har den breda demokratiska bas som �r n�dv�ndig f�r att �terinf�ra etnisk harmoni och att hj�lpa landet ur den ekonomiska svacka som det nu befinner sig i .
frankrike accepterar av samma sk�l alla de tarvligheter som dess beskyddare i den ivorianska statens ledning g�r sig skyldiga till , bara de i geng�ld skyddar de franska intressena .
m�nskliga r�ttigheter
antalet politiska f�ngar f�refaller ha �kat fr�n 1 500 till 3 000 helt nyligen , och m�nga av dem tvingas att utf�ra straffarbete och �r utsatta f�r grymma former av tortyr .
problemet �r naturligtvis vad vi nu , som europeiska unionen , kan g�ra ?
herr talman ! jag har i m�nga �r haft en affisch p� v�ggen i mitt kontor av aung san suu kyi n�r hon tilldelades sacharovpriset av detta parlament .
ett stort antal av dem har arresterats eller trakasseras och f�rs�k har gjorts att st�nga deras huvudkvarter i burma .
n�r allt kommer omkring har v�st spelat en viss roll i vietnam .
det kr�vs s�ledes att europeiska unionen b�rjar inta en beslutsam attityd i f�rh�llande till vietnam och st�ller fr�gan om r�ttsstatsprinciper , och inte bara - jag upprepar det - fr�gan om de m�nskliga r�ttigheterna , som man kan notera har f�rb�ttrats n�got .
jag vill bara be om att man hanterar denna sak med f�rsiktighet , och jag hoppas att ni urs�ktar att jag missbrukar talartiden som g�ller vietnam .
kriget mellan de tv� l�nderna har inte lett till n�gon permanent f�rbittring .
president clinton skulle g�ra gott i att ta upp detta i hanoi under sitt bes�k .
vietnam har sedan dess till�mpat en utrikespolitik med �ppna d�rrar . tack vare den upptar landet den plats den �r v�rd i v�ra internationella f�rh�llanden .
vi vet ju vad det handlar om .
detta �r naturligtvis en klen tr�st f�r de som lever med smutsigt vatten som rinner genom deras hus och som kan komma att st�llas inf�r enorma ekonomiska f�rluster .
detta �r otvivelaktigt sant .
det �r inte r�ttvist att m�nniskor skall beh�va uppleva tragedier av denna proportion och sedan konfronteras med en mycket os�ker framtid eftersom klimatf�r�ndringarna redan sker , och de problem som de har upplevt under de senaste tv� veckorna �terkommer s�kerligen , om inte under n�sta �r , s� s�kert under de kommande �ren .
d�rf�r �r det dessa industrier som m�ste anstr�nga sig mest f�r att minska utsl�ppen .
tack s� mycket , herr kommission�r .
och nu �r det tanken att vi skall r�sta om en s� pass viktig text med ett deltagande som uppskattats till 171 ledam�ter !
jag respekterar de kommentarer ni har gjort och kan f�rs�kra er om att de kommer att bli inf�rda i protokollet .
f�r eu har principen om en fri tj�nstesektor st�rre betydelse �n r�tten till h�lsa och v�rd , och den underminerar d�rigenom metodiskt och systematiskt det offentliga h�lso- och sjukv�rdssystemet , s�rskilt inom omr�det f�r v�rd , med det anst�tliga gynnandet av de privata f�rs�kringsformerna som ett " n�dv�ndigt " komplement eller t.o.m. substitut f�r den offentliga sociala tryggheten .
trots korrekta �verv�ganden om vilken niv� vi har uppn�tt med de befintliga systemen , som syftar till att ge varje medborgare en h�g skyddsniv� oberoende av egna resurser och individuella risker ; trots en betoning av riskerna med �verflyttningar mellan offentliga och privata system ; trots en beskrivning av att deras andel av de totala utgifterna �kar och de oj�mlika f�rh�llanden som uppst�r d�rvidlag - trots allt detta �r alla konkreta f�rslag i resolutionen inget annat �n en uppmuntran till att gemenskapen skall p�skynda utvecklingen av privata f�rs�kringssystem .
alla tvingas att endast visa solidaritet med sig sj�lva , och att �gna sig �t alla m�jliga on�diga penningaff�rer .
kapitalbas i kreditinstitut ( forts . )
bara p� s� vis kan man ju skapa likadana konkurrensvillkor .
men det faktum att det l�ggs fram , i likhet med kommissionens nya initiativ , �r d�remot n�got som kan verka f�rv�nande .
vi s�ger " ja " till en starkare inriktning av kapitalt�ckningen betr�ffande kreditrisker p� det ekonomiska riskinneh�llet och till en vidareutveckling av f�reskrifterna om egna medel .
. ( es ) herr talman ! f�r det f�rsta skulle jag vilja uppm�rksamma att kommissionen med tillfredsst�llelse ser att villiers bet�nkande inte bara p�verkar utv�rderingen av kapitalbasdirektivet utan ocks� den aktuella �versynen av �ndringarna i f�rordningarna om utj�mning av kapital .
vi b�r st�dja dessa m�l med hj�lp av v�l �vert�nkta , s�kra regler som garanterar v�ra marknaders och v�ra institutioners s�kerhet .
jag f�rklarar debatten avslutad .
med tanke p� att vi h�r i parlamentet inom kort m�ste b�rja arbeta med betydande f�r�ndringar av stadgan f�r europeiska ombudsmannen , vilka fortfarande diskuteras i utskottet f�r konstitutionella fr�gor , och vars bet�nkande ocks� har anf�rtrotts mig och handlar om utvidgningen av unders�kningsbefogenheter f�r ombudsmannen , reserverar vi den kvalitativa och kompletta revideringen av texten i respektive stadga till denna tidpunkt .
ombudsmannens kansli bidrar sannerligen till att ge oss uppr�ttelse f�r denna brist p� demokrati .
jag f�rklarar debatten avslutad .
det �r hennes uttryckliga �sikt som jag vill f�sta uppm�rksamhet vid n�r jag talar ikv�ll .
herr talman ! b�sch har lagt fram ett utm�rkt bet�nkande , som han b�r tackas f�r , vilket ocks� hautala har gjort f�r utskottet f�r r�ttsliga fr�gor .
f�redraganden f�r europaparlamentets utskott f�r framst�llningar konstaterar i motiveringarna till bet�nkandet att de principer som ledde till de rekommendationer som ombudsmannen formulerat visat sig �verensst�mma med europaparlamentets , n�mligen korrekthet , �ppenhet och en �nskan om att inge f�rtroende .
ombudsmannens initiativ och rekommendationer v�lkomnas d�rf�r varmt , liksom kommissionens beslut att f�lja dem .
vi kunde inst�mma vem som helst i landet inf�r ombudsmannens utskott , och det s�rskilda utskottsf�rfarandet , vilket jag kommer att diskutera p� tv� minuter , �r n�got som vi kan l�ra av .
europeiska unionen har en kort historia till skillnad fr�n medlemsstaterna som har ett l�ngt f�rflutet . och d�rf�r m�ste den skapa f�rhoppningar om n�got nytt .
slutligen kan kommissionen naturligtvis sj�lv g�ra egna �taganden .
justering av protokollet fr�n f�reg�ende sammantr�de
ett s�tt att vinna omr�stningar �r att vara n�rvarande n�r dina motst�ndare inte �r det .
. ( it ) jag r�stade f�r villiers bet�nkande om kapitalbasen i kreditinstitut , eftersom direktiv 89 / 299 / eeg som antogs f�r att reglera detta omr�de f�r hela elva �r sedan m�ste uppdateras och kompletteras .
vi st�der kravet p� att man m�ste hitta en l�sning p� den konflikt mellan usa och eu som �r en f�ljd av den diskriminerande gramm-leach-bliley-lagstiftningen .
jag tackar den bayerska och den tyska inrikesministern liksom �sterrikes f�rra inrikesminister schl�gel , som gemensamt m�jliggjorde detta vid m�tet i tammerfors .
naturligtvis b�r �ven de l�nder prioriteras med vilka europeiska unionen f�r f�rhandlingar om anslutning .
n�r en person suttit h�ktad i 110 dagar utan r�tteg�ng m�ste han friges och kan aldrig mer �talas f�r samma brott .
jag tar ett exempel . posselt skriver : genomf�rande av kurser f�r nationella poliser p� basis av gemensamma normer .
karamanou sade alldeles nyss att han var glad �ver att europaparlamentet kommer att f� en r�dgivande roll . bara h�romdagen r�stade den socialistiska gruppen emot , f�r i europols styrelse fanns det parlamentsledam�ter med r�str�tt .
om en siare p� den tiden hade varnat f�r att det skulle sluta med att den lokala kvarterspolisen visslar " ode till gl�djen " och f�rs�ker lista ut hur man skall till�mpa det europeiska tillv�gag�ngss�ttet p� polisarbetet i kurran skulle ingen i storbritannien n�gonsin ha trott honom .
parlamentet kan vara stolt �ver att f�rslaget att inr�tta denna akademi f�ddes h�r och vi �r tacksamma f�r att det portugisiska ordf�randeskapet tog upp f�rslaget och f�r att kommissionen och r�det st�der det .
vi ser att polisen i det ena landet reagerar helt annorlunda p� samma situation �n i det andra landet .
framf�r allt vill jag understryka att enligt dem som till exempel alltid har f�rsvarat en n�rpolis , som n�r det g�ller f�renade kungariket , skulle jag vilja gratulera till att detta begrepp med brittiskt ursprung f�r allt st�rre st�d hos en rad l�nder i det s� kallade kontinentala europa .
som parlamentsledam�ter ber�rs vi sj�lva mycket ofta av kriminalitet .
vidare skulle akademins organisation vara flexibel och r�rlig , utbildningen skall kunna �ga rum i varje enskilt fall vid den mest kvalificerade nationella h�gskolan .
jag har arbetat med dessa fr�gor i �ver sex �r och haft flera betydande framg�ngar med att h�mta tillbaka bortf�rda barn , till stor del tack vare europaparlamentets st�d och resurser .
emellertid beklagar vi att till�mpningsomr�det f�r denna f�rordning begr�nsas , att den inte omfattar ogifta par , d�r barn har f�tts utanf�r �ktenskap , vilka d�rigenom inte f�r sina r�ttigheter erk�nda och till�mpade inom gemenskapsramen .
detta �r en uppgift f�r framtiden .
men jag har �nnu fler inv�ndningar mot att man angriper juridiska svagheter och prejudicerande effekter , vilket leder till att ett samh�llsproblem l�mnas utan l�sning f�r �versk�dlig framtid .
herr talman ! jag tvivlar inte ett �gonblick p� kommission�r vitorinos engagemang i denna fr�ga .
kommissionen anser att det g�llande f�rdraget om europeiska unionen g�r det m�jligt att ta h�nsyn till idrottens egna s�rdrag i allm�nhet , och dess sociala funktion i synnerhet .
jag vet hur engagerad och besluten den �r att g�ra detta och jag vet naturligtvis ocks� att idrott och s�rskilt fotboll handlar om stora aff�rer och inte kan v�ntas vara undantagen fr�n vanliga regler f�r f�retagsverksamhet .
europaparlamentet har ofta gett utryck f�r oro i dopningsfr�gan och kr�vt effektivare mot�tg�rder .
d�rmed har vi behandlat denna punkt .
detta f�rslag �r speciellt h�rt och f�rargligt f�r irland .
det vi m�ste klara ut i dag �r att f�renade kungariket f�resl�r det den g�r fullt medveten om att den m�ste samr�da med europeiska unionen och fullt medveten om att det finns gemenskapslagstiftning som den m�ste f�lja .
jag hoppas verkligen att detta kommer att bli ett av resultaten av detta .
jag lyssnade p� mccartin tidigare och det �r uppenbart att han har missuppfattat detta fullst�ndigt .
en lokal �kare i danmark eller i f�renade kungariket f�r valuta f�r sina pengar 365 dagar om �ret , men en utl�ndsk �kare fr�n n�gon annan medlemsstat som k�r in i landet - kanske f�r att stanna en eller tv� eller tio eller till och med hundra dagar - f�r det inte .
tyv�rr har ett nytt v�ldsbudskap riktats mot v�ra demokratier , med det s�rskilt f�rhatliga mordet p� ernest lluch .
ni vet att vi har en fullsp�ckad f�redragningslista , och med st�d av de befogenheter som arbetsordningen ger mig f�r att se till att kammarens arbete fungerar v�l , har jag s�ledes fattat detta beslut .
efter intensiva f�rhandlingar , b�de p� teknisk niv� och ministerniv� , p� grundval av f�rslag till beslut med ca 500 parenteser , blev det inte m�jligt att sluta ett helt�ckande avtal om de viktigaste politiska sakfr�gorna .
det framgick till sist , emellertid , att eftergifterna fr�n andra parter om " komplementaritet " , efterlevnad och kyotomekanismerna var otillr�ckliga f�r att kompensera f�rsvagningen av m�len f�r utsl�ppsminskningen , som hade blivit resultatet om f�rslagen om " kols�nkor " hade godk�nts .
det var , p� s�tt och vis , en v�ntad olycka - som titanic och isberget .
hos oss tilltar utsl�ppen med koldioxid , det vet vi och det har vi tillr�ckligt ofta diskuterat h�r .
fru talman ! konferensen om v�rldens klimat har misslyckats , men trots det kan man notera verkliga framg�ngar .
lyckligtvis var 14 av de 15 milj�ministrarna �verens om detta .
enligt den andra uppfattningen har europeiska unionen misslyckats eftersom tysklands och frankrikes " gr�na " milj�ministrar inte var beredda att gl�mma kyoto .
detta kyotoprotokoll f�r inte under n�gra omst�ndigheter urvattnas .
om det g�r att n� ett avtal med f�renta staterna om ett l�gre faktiskt genomf�rande i eget land , s� �r det alltid b�ttre �n inget avtal �ver huvud taget .
l�t oss trots allt avsluta med en hoppfull notering .
vi har sj�lva alltid sagt att inget avtal �r b�ttre �n ett d�ligt avtal , men det betyder inte att vi kan g�ra v�r egen politiska �nskelista till en m�ttstock f�r ett bra avtal .
fru talman , �rade ledam�ter ! jag vill som ordf�rande f�r europaparlamentets delegation f�r cop6 , b�rja med att gratulera till det utm�rkta f�rh�llande som kommissionen och parlamentet har haft under denna vecka .
nu �r det l�ge att best�mma oss f�r att vi inte skall kunna misslyckas en g�ng till .
vi inledde diskussioner om vad vi tidigare hade bed�mt vara stora kryph�l , eller m�jliga stora kryph�l .
vi har n�jet att v�lkomna minister hubert v�drine .
n�r det g�ller fr�gan om kvalificerad majoritet har arbetet framskridit . med vissa medlemmars anstr�ngningar , om dessa bekr�ftas , skulle ett trettiotal best�mmelser kunna omfattas av omr�stningar med kvalificerad majoritet .
en str�mning �r m�jlig att uppfatta - jag s�ger det med f�rsiktighet eftersom flera medlemsstater kanske �nnu inte kommit fram till en slutlig st�ndpunkt i fr�gan - men det g�r att uppfatta en str�mning till f�rm�n f�r enkel viktning , �ven om det naturligtvis �terst�r att sl� fast omfattning och exakta villkor .
de har t.o.m. planerat att toppm�tet skall kunna p�g� �ven under s�ndagen om detta visar sig vara n�dv�ndigt .
m�tet i nice blir ett tillf�lle till att diskutera unionens institutionella reform med alla kandidatl�nder , och mer generellt europas framtidsutsikter .
i den andan - i lissabons efterf�ljd - har det franska ordf�randeskapet bl.a. prioriterat ett antagande av den sociala dagordningen .
inf�r europeiska r�dets toppm�te f�rbereds slutligen en f�rklaring om idrottens ekonomiska , sociala och kulturella s�rdrag samt sociala funktioner i europa .
( appl�der ) naturligtvis anser medlemsstaterna att det �r politiskt sv�rt att avst� fr�n vetor�tten p� k�nsliga omr�den som socialpolitik , asyl- och invandringspolitik , gemensam handelspolitik , sammanh�llning och skatter �ven n�r man bara talar om de tekniska f�r�ndringar som erfordras f�r att f� den inre marknaden att fungera .
vi anser ocks� att ni betr�ffande fr�gor , d�r vi �nnu inte uppn�tt n�got majoritetsbeslut , i f�rdraget redan kan skriva in att man genom ett enh�lligt beslut , med iakttagande av vissa tidsfrister , kan �verg� till majoritetsbeslut , ty om man skriver det s� i f�rdragen , beh�ver man inte varje g�ng g�ra en revidering av f�rdragen med ett utdraget ratificeringsf�rfarande .
f�r det andra anser vi att man inte b�r g� fram�t bara n�r det g�ller kvalificerade majoriteter , utan att det alltid m�ste vara medbeslutande i lagstiftnings�renden .
min v�djan till er , herr r�dsordf�rande , �r att ni l�gger fram ett dokument f�r oss i detta parlament som �r tillr�ckligt bra f�r att godk�nnas av oss , och som ocks� �r ett dokument som lever upp till den stora historiska utmaning vi st�r inf�r i europa .
jag s�ger att om vi kompromissar och s�tter ribban f�r l�gt , kommer vi att v�gra ta detta p� allvar , och det g�r vi f�r europas b�sta och med gott samvete .
detta skulle vara ett ytterst betydelsefullt st�llningstagande av parlamentet , vilken vi kan r�sta om i morgon .
troligt �r att man kommer att fatta beslut om �tg�rder under den sista natten , beslut som v�ra nationella parlament inte uttryckligen har diskuterat , och som man sedan kommer att be dem ratificera i den obligatoriska kompromissens namn .
det finns fortfarande 65 best�mmelser kvar med enh�llighet i amsterdamf�rdraget .
i demokratier �r det tv�rtom .
det �r emellertid inget svar p� den inst�llsamhet i beslutsprocessen som fortfarande r�der h�r inom europeiska unionen .
alla , eller n�stan alla , har sagt det f�re mig : vi vill att stadgan skall omn�mnas i artikel 6.2. underskatta inte parlamentets beslutsamhet att uppn� detta .
dess r�st skulle bli starkare , och de ministrar som f�rsvarar jordbruket , det jordbruk som gynnar en h�llbar utveckling , skulle ocks� f� en starkare r�st i r�det om de kunde st�dja sig p� beslut som fattats h�r i enlighet med medbeslutandef�rfarandet .
herr talman ! jag deltog aktivt i den danska folkr�relsen mot maastrichtf�rdraget 1992 .
herr talman , herr r�dsordf�rande , herr kommissionsordf�rande ! den lettiska presidenten har i dag vid ett samtal i kammaren f�rebr�ende sagt - med adress till oss : vi g�r v�ra heml�xor !
jag vill p�peka att befolkningen ser sig f�retr�dd av europaparlamentet , och det m�ste komma till uttryck i europaparlamentet !
herr talman ! till och med i paris r�der delade uppfattningar om nice .
stadgan f�rtj�nar inte att bli h�ngande i tomma luften utan tydlig status .
sedan beh�ver man inte t�nka s� l�ngt f�r att inse att antalet 700 parlamentsledam�ter inte l�ngre kan g�lla f�r ett europa med tjugosju eller tjugo�tta nationer , utan att de mindre l�nderna f�r uppleva en minskning som jag anser vara or�ttvis .
herr talman , herr r�dsordf�rande , herr kommissionsordf�rande ! omedelbart efter m�tet i nice n�rmar sig den tidpunkt d� europaparlamentet uppmanas svara p� tv� historiska fr�gor , den ena g�ller europeiska unionens framtid och den andra parlamentets egen politiska trov�rdighet .
detta �r naturligtvis viktigt och jag �r �verraskad att ingen annan har n�mnt det , eftersom det tagit upp s� mycket av v�r tid i utskottet .
efter president chiracs tal h�r i juli m�nad vet vi att �tminstone tre stora fr�gor kommer att klarg�ras , n�mligen en f�renkling av f�rdragen ; befogenheterna p� europeisk , nationell och regional niv� , n�got jag skulle kalla staternas r�ttigheter enligt ett amerikanskt uttryck - artikel 10 i den amerikanska konstitutionen - och f�r det tredje j�mvikten mellan institutionerna . men i den fr�gan �r det kanske de nationella parlamentens roll som b�r �verv�gas i f�rsta hand , dvs. hur v�r institution skall f�rvaltas i framtiden .
det �r inget att vara r�dd f�r .
n�r det g�ller det ut�kade bruket av kvalificerad majoritet inst�mmer vi i att om vi inte tar vissa steg i riktning mot ut�kning kommer vi att f� v�ldigt m�nga problem .
det som h�nt vike freiberga �r belysande f�r hur central- och �steuropas folk b�r sina sv�righeter med j�mnmod .
som kollega ber�s sade �r det naturligtvis en oh�llbar �tskillnad att vi � ena sidan har medbeslutander�tt i konsumentfr�gor och samtidigt endast yttrander�tt i jordbruksfr�gor .
n�r vi lyssnar p� bonde , s� �r balkan hans slutliga ideal .
denna g�ng �r det visserligen , paradoxalt nog , det samf�rst�nd som kan sk�njas som ger m�nga av oss politisk huvudv�rk .
herr talman ! vi fr�n forza italia och ppe tror p� detta och kommer att st� vid er sida under byggandet av medborgarnas europa .
n�r vi v�l n�dde ett samf�rst�nd om den h�r texten , som f�r �vrigt �r en bra text , mycket v�l f�rberedd av konventet , en text som �r l�tt att l�sa , som har stil , d� s�ger vissa l�nder : den m�ste integreras i artikel 6 .
n�r vi utvecklade id�n att vi i framtiden kommer att ha ett intresse av att kommissionen inte blir alltf�r stor , f�r att den skall kunna f�rbli effektiv och beh�lla all sin kapacitet , framf�r allt sin initiativmakt , visade vi att ocks� vi var beredda att g�ra den uppoffringen .
jag tackar er �n en g�ng - tillsammans kommer vi att hitta den l�sningen .
jag f�rklarar debatten avslutad .
herr talman ! jag skulle vara tacksam om ni rapporterade till kammaren om de fr�gor som jag har tagit upp .
herr talman ! jag k�nde inte till den incidenten .
jag kan meddela er att fontaine , enligt vad jag erfarit och vilket jag inst�mmer i f�r presidiets r�kning , beklagar den h�r allvarliga incidenten mycket djupt .
herr talman ! i g�r intr�ffade n�gonting enormt allvarligt i italien .
detta utm�rkta initiativ f�rnyades i �r , och det andra forumet kommer att h�llas den 12 och 13 december i paris , dvs. under europaparlamentets sammantr�desdagar i strasbourg .
herr gorostiaga ! jag fr�ntar er ordet .
h�r inst�mmer vi ocks� i att rangordningen �r riktig .
herr f�rsvarsminister ! vi gl�der oss �t detta .
det finns �ven m�nga andra saker att ta upp . genom att v�nda mig till r�dets f�retr�dare skulle jag vilja tala om f�r dem att europaparlamentets vilja �r att vi skall f�rv�rva denna s�kerhets- och f�rsvarskultur , som vi inte har n�gon vana vid , och vi �nskar att toppm�tet i nice blir en odelad framg�ng .
de institutionella aspekterna �r ocks� mycket viktiga , eftersom de g�r att unionen kan f�rutse , besluta och agera , dvs. s�kerst�lla den politiska kontrollen och den strategiska ledningen i en krishanteringsoperation .
som brok �nskar i sitt bet�nkande , kommer r�det att f�rfoga �ver register som sammanfattar alla f�rbindelser mellan unionen och vart och ett av partnerl�nderna , f�r att kunna dra st�rre nytta av unionens sammantagna utgifter , �ka deras effektivitet och b�ttre f�rbereda sina debatter i fr�ga om externa �tg�rder .
i det h�r sammanhanget var det toppm�te som nyligen h�lls i zagreb mycket viktigt .
ordf�randeskapet har �gnat sig �t att utveckla unionens f�rbindelser med andra stora regionala enheter och m�nga asiatiska m�ten : det tredje asem-toppm�tet , toppm�tet med japan och med kina .
jag skulle vilja kunna s�ga att v�ra p�tryckningar och �tg�rder p�verkar den nuvarande situationen . tyv�rr finns det en sorts motst�nd och autonomi i den afghanska situationen inf�r alla dessa insatser .
dels en kapacitetskatalog , dvs. ett dokument p� 300 sidor som noggrant identifierar den milit�ra kapacitet som unionen anser n�dv�ndig f�r att fullg�ra samtliga petersberguppdrag .
det �r s�ledes en ny dynamik som har satts ig�ng , p� grundval av en politisk viljehandling fr�n medlemsstaternas sida .
. ( en ) jag kanske kan b�rja med att kommentera vad min hederv�rde v�n hume just har sagt .
precis som ministrarna p�pekat i sina utm�rkta tal , har vi under de senaste veckorna bevittnat en viktig utveckling n�r det g�ller att st�rka europas bidrag till sin egen s�kerhet .
utmaningen f�r oss nu �r att h�lla fast vid denna strategi , se till att vi kan f� denna strategi att fungera och se till att , genom att h�lla d�rren �ppen f�r n�rmare f�rbindelser med den europeiska familjen , vi kan hj�lpa dessa l�nder att genomf�ra de ekonomiska och politiska f�r�ndringar och reformer som kr�vs f�r att s�kra deras stabilitet och l�ngsiktiga v�lst�nd .
n�r det g�ller tillhandah�llandet av bist�nd , har kommissionen fr�mst genom sitt kontor f�r humanit�rt bist�nd , echo , gjort en rad specifika interventioner i �r som syftar till att lindra b�da effekterna av den katastrofala torkan i landet genom att st�dja - genom tillhandah�llande av medel f�r livsmedelss�kerhet och utrustning inf�r vintern - de befolkningsgrupper som f�rdrivits p.g.a. striderna i den nord�stra delen av landet .
nu g�ller det ocks� att med detta som utg�ngspunkt forma en effektiv , rationell europeisk enhet som skall st� under entydig ledning .
herr talman , herr r�dsordf�rande ! ofta tar det mycket l�ng tid innan synliga resultat kan sk�njas n�r fr�gor behandlas p� europeisk niv� .
det inneb�r att det m�ste finnas strukturer f�r oss parlamentariker f�r att vi skall kunna f� information om besluten , kunna debattera , delta och utkr�va ansvar .
den f�rsta �r europaparlamentets roll , vilket ett flertal kolleger ocks� har n�mnt .
jag kan tala om att palestiniernas f�rv�ntningar p� europa �r �verv�ldigande .
som en organisation med soldatm�drar h�vdar : vi har inte h�mtat hem v�ra barn fr�n libanon f�r att de skall d� f�r bos�ttningarna .
konflikten i mellan�stern skulle d�rf�r kunna bli en sorts bekr�ftelse p� effektiviteten i den europeiska mellan�sternpolitiken .
herr minister , jag vill s�rskilt tacka f�r att ni var i utskottet och att ni �r h�r i dag .
d� kunde de �vriga eu-l�nderna h�lla sig till traditionell fredsbevarande verksamhet .
den kan bara �tervinna sin trov�rdighet om den har en civil inriktning som f�rsta princip , om den bedriver en effektiv f�rebyggande politik med de instrument som st�r till f�rfogande , och �ven utrustar dessa ekonomiskt p� ett trov�rdigt sett .
mot den fienden riktar sig er gusp .
f�r det andra : nato b�r stegvis uppl�sas och inte utvidgas �sterut .
jag kan inte uttrycka hur glad jag �r att uppt�cka att brok hela tiden har varit en farlig revolution�r !
det vi nu �gnar oss �t �r att p� alla s�tt st�rka f�ruts�ttningarna f�r frihet och fred i europa .
jag tror att om vi kunde f�rst� detta klart och tydligt , skulle kanske mycket av oron f�rsvinna .
det �r n�dv�ndigt att garantera en demokratisk kontroll av hela denna process .
precis som min fine gael-kollega , doyle , inser jag att detta inte �r detsamma som skapandet av en europeisk arm� , och innan det blir ett alltf�r h�gljutt klagande i mitt hemland , vilket det kommer att bli , mot irlands deltagande , vill jag p�peka att deltagandet �r frivilligt och att det bed�ms fr�n fall till fall .
alla politiska och diplomatiska anstr�ngningar och ekonomiska p�tryckningar kunde inte f�rhindra ett v�ldsutbrott i europas hj�rta och en oacceptabel utmaning av alla europeiska v�rderingar .
jag kan f�r �vrigt konstatera att det i r�dets alla st�ndpunkter inte finns och inte kommer att finnas ett budget�rt �tagande f�r europeiska unionen att finansiera n�gon som helst milit�r verksamhet .
a5-0326 / 2000 av harbour , f�r utskottet f�r r�ttsliga fr�gor och den inre marknaden , om kommissionens vitbok om reformen av kommissionen ( aspekter som ber�r utskottet f�r r�ttsliga fr�gor och den inre marknaden ) ( kom ( 2000 ) 200 - c5-0446 / 2000 - 2000 / 2216 ( cos ) )
d�rf�r �r vi m�na om att den inte skall beh�va lida , men det �r mycket viktigt f�r oss att all personal verkligen �r delaktig i hela denna moderniseringsprocess .
en �rlig utv�rdering av organisationens utveckling och merkostnaderna f�r reformen kr�ver en samordning i b�rjan av varje budget�r .
dessutom �r det helt ologiskt att endast r�det skall kunna �ndra p� de finansiella best�mmelserna , och vi upprepar v�r beg�ran om f�rlikning p� den punkten .
och vi har ocks� varit enh�lliga i att konstatera att en stor del av de brister och oegentligheter som man klagade p� under godk�nnandet av f�rvaltningen �r 1996 berodde p� det faktum att tidigare kommissioner varken lyckades modernisera sina f�rvaltnings- och kontrollsystem eller i sin helhet till�mpa g�llande regler .
ett bevis p� denna svaghet �r det oerh�rt begr�nsade antalet avslag p� godk�nnanden , p� tillst�nd , av kommissionen .
det jag tyckte var mycket intressant , var att diskussionerna visade hur syssels�ttnings- och organisationspraxisen inom den privata och offentliga sektorn faktiskt b�rjar bli allt mer lika .
ledarskap fr�n toppen kommer att bli n�dv�ndigt .
det �r till sist ocks� dags att intressera sig f�r unionens externa representation .
d�rf�r fr�gar vi kommission�ren : kan kommissionen garantera en �verg�ngsperiod som i tiden verkligen �r begr�nsad ?
det gl�der mig att det verkar som om kommissionens f�rslag verkar vara f�renligt med den st�ndpunkt som vi skall anta i morgon .
cheferna f�r enheterna och organen b�r ha en viss r�relsefrihet betr�ffande administrationen .
h�r ser vi fortfarande att det finns en del att ta igen , och vi hoppas p� att kommissionen v�gar vara �ppnare .
herr talman ! i sitt brev till romarna uppmanar aposteln paulus sina l�sare att omdana sig genom att f�rnya sitt t�nkande .
herr talman , �rade ledam�ter ! f�rden mot de nya europeiska institutionerna forts�tter i och med f�rslaget till en reformering av kommissionen : jag s�ger " nya " eftersom de kommer att f�r�ndras j�mf�rt med tidigare till f�ljd av de problem som uppstod under den f�rra ledningen och p� grundval av den l�nga , m�ngfacetterade och ofta komplicerade rapporten fr�n de oberoende experterna .
som ni kanske f�rv�ntade er , st�der vi �ndringsf�rslag 1- 6 , som ingetts av pse-gruppen .
n�r det r�r utvidgningen , s�ger lamassoure att kommissionen , n�r det g�ller anslutningsprocessen , f�rv�ntas l�gga fram en helt�ckande strategi som �terspeglar unionens intresse av dess politiska tidtabell - inte bara en bed�mning med h�nsyn till varje enskilt ans�karlands l�mplighet .
med beaktande av detta uppmuntrar vi kommissionen och kinnock att fullf�lja sitt reformarbete .
herr talman ! kommissionens avg�ng v�ren 1999 utgjorde i sj�lva verket finalen f�r ett l�ngt mer djupg�ende problem hos europeiska kommissionen : otydligt definierade arbetsstrukturer som resulterade i en brist p� politiskt ansvar , splittrade politiska prioriteringar och otillr�ckliga resultat .
detta kan inte uppn�s med en f�r stor fokusering p� ordet " intern " i reformerna .
utrikesfr�gor �r viktiga och intressanta f�r europaparlamentet , och eftersom jag sj�lv haft ett livsl�ngt intresse f�r s�dana fr�gor , tror jag att detta �r en korrekt f�rklaring .
man betonar ansvaret f�r dem som tar emot uppgifter om m�jliga oegentligheter att agera snabbt , seri�st och effektivt .
jag �r �vertygad om att kammaren kommer att ge er m�jlighet att utbreda er mer vid ett annat tillf�lle , med tanke p� att denna reform inte kommer att vara avslutad i och med den f�rsta omr�stningen i morgon .
allts� , �n en g�ng , m�let �r �ppenhet , och jag tror att vi kommer att uppn� detta m�l .
d� gl�mmer man ofta bort att vi ocks� lever i ett demokratiskt system d�r vi har regler om medbeslutande , och det �r bra .
kommissionen bibeh�ller , �ven om det �r sant att det sker p� ett nyanserat s�tt , en uppdelning mellan det politiska ansvaret och den verkst�llande befogenheten , som vi av tidigare erfarenhet f�rutser att den inte kommer att vara s�rskilt operativ .
( talmannen uppfordrade talaren att avsluta sitt inl�gg . ) herr talman , jag skall avsluta med att s�ga att vi kommer att godk�nna tv� �ndringsf�rslag och avsl� tre , som vi redan diskuterat i kommissionen .
det �r ett mycket bra initiativ av sauquillo att ocks� ta med delen om utl�ndska f�rbindelser i samband med den interna reformen och d�rmed ocks� f�ra upp detta p� f�redragningslistan .
fattigdomen och n�den beror inte bara p� ekonomisk underutveckling och utvecklingssv�righeter utan �r ofta resultat av att de starka angriper och utnyttjar de svaga , av de dugligas egoism gentemot de utslagnas svaghet .
vi b�r slutligen f�rst� att kommission�r pattens f�rslag om att en styrelse best�ende av ledam�ter fr�n kommissionen , med kommission�r nielson som verkst�llande direkt�r skall vara ansvarig f�r bist�ndet , �r ett ogenomf�rbart p�fund som l�nats ur managementlitteraturen och i grunden �r of�renligt med kommissionens kollegiala struktur .
v�rt utskott delade f�redragandens uppfattning att det �r kommission�ren ansvarig f�r bist�nd som b�de skall formulera och verkst�lla politiken inom detta omr�de , �ven om den skall samordnas med �vriga politikomr�den som handlar om utrikes verksamhet .
h�r har �terigen budgetmyndighetens f�rst�else spelat en avg�rande roll f�r finansieringen av denna omfattande omorganisation av eu : s tj�nst f�r yttre f�rbindelser .
( sammantr�det avbr�ts kl . 00.30. )
fr�mst i frankrike s�ger somliga till mig att vi m�ste vidta kraftfulla nationella �tg�rder f�r att skydda den franska kusten , och en del f�resl�r rentav att vi skall inf�ra franska kustvakter .
. ( en ) fru talman ! jag anser att det inte r�der n�gon tvekan om att kommissionen i likhet med det franska ordf�randeskapet anser att fr�gan om sj�s�kerhet och milj�skydd �r ytterst viktig .
jag vill avsluta med att tacka herr gayssot , ordf�rande i ministerr�det ( transport ) , f�r hans stimulerande synpunkter .
vi �r alla �verens om det , men vi m�ste hitta en metod med vilken denna prioriterade �tg�rd kan genomf�ras och �nnu har vi inte n�tt en �verenskommelse mellan de tre institutionerna om det .
som watts redan har f�rklarat s� har europaparlamentet p� flera punkter en str�ngare uppfattning �n vad r�det tycks ha .
utskottet har �ven haft m�ten med ber�rda sektorer och m�nga kontakter har tagits med det franska ordf�randeskapet i syfte att kunna komma fram till en text som alla parter kan samtycka till och som kan godk�nnas snabbt av de tv� lagstiftande institutionerna : r�det och europaparlamentet .
�ven om industriellt och radioaktivt utsl�pp forts�tter fr�n en rad k�llor anses nu allm�nt praxis med direkt dumpning med lite tanke p� framtiden vara oacceptabelt .
allm�nheten har dessutom r�tt att f� veta vilka f�rberedelser som har gjorts , vilken typ av material som utg�r en fara och vilka f�ljder som kan f�rv�ntas .
jag �r �vertygad om att detta p� sikt m�ste leda till att vi inr�ttar en europeisk kustbevakning .
jag kommer att st�dja detta bet�nkande och kommissionens �ndringar , men jag uppmanar ledam�terna att �ven st�dja �ndringarna fr�n utskottet f�r milj� r�rande sociala normer .
mindre gl�djande , och det p�mindes vi just om , �r att staterna i europeiska unionen i det f�rg�ngna sannerligen inte har sk�rdat n�gra lagrar n�r det g�ller s�kerhet p� fartyg .
var sn�ll och hj�lp till s� att kommissionen h�r ger en tydlig signal .
var och en som jobbar inom den sektorn har ett tungt ansvar .
herr talman , fru kommission�r , herr tj�nstg�rande r�dsordf�rande ! de senaste m�nadernas katastrofer har kastat ljus �ver det otillr�ckliga regelverket , bristerna vad avser kontrollsystem och m�nskliga och finansiella resurser .
f�r n�gra veckor sedan drabbades v�stra frankrike av en ny ekologisk katastrof , d� kemikaliefartyget ievoli sun havererade . och det �r f�rst i dag som europaparlamentet finner anledning att uttala sig om en �kad sj�s�kerhet .
helt riktigt pekar f�redraganden p� att det skick som en tankb�t befinner sig i s�ger mer �n dess �lder .
herr talman ! jag begr�nsar mig till att kommentera och framf�ra den �sikt som majoriteten av den socialistiska gruppen hyser om ett av �ndringsf�rslagen , det f�rslag som �ndrar det direktiv som reglerar inspektionsmyndigheterna .
vi vill inte ha dem i v�ra farvatten och inte i v�ra hamnar .
jag skall nu koncentrera mig p� tv� �renden : hamnstatskontroll och utfasning av oljefartyg med enkelskrov .
om vi skall bli trov�rdiga m�ste vi handla snabbt och avbryta den politiska retorik som inte leder till n�got konkret .
alla k�nner vid det h�r laget varandras inst�llning och �ven av den anledningen beh�ver vi f�reta omr�stningen i dag !
det finns emellertid �nnu mycket att g�ra inom denna sektor .
r�ttvisan vet att vara skoningsl�s mot fattiga som inte kan betala en avgift eller b�ter , och g�r s� l�ngt som till att beslagta deras ynka �godelar .
jag anser d�rf�r att det �terst�r oerh�rt mycket att g�ra p� detta omr�de .
det �r d�rf�r viktigt att sl� fast vissa politiska och kulturella grundf�ruts�ttningar : vi m�ste sluta t�nka i termer av katastrofer och i st�llet b�rja koncentrera oss p� f�rebyggande arbete .
s�kerhetsproblemet hos transporterna m�ste l�sas genom rationella sanktioner av lag�vertr�darna , sanktioner som medf�r kostnader f�rdelade �ver sektorn p� global niv� , s� att vi inte skadar den europeiska sektorn �nnu mer .
n�r vi g�r detta m�ste vi alltid komma ih�g att dubbelskrov eller till och med tredubbla skrov inte med absolut s�kerhet garanterar att olyckor inte kommer att �ga rum i framtiden .
till herr jarzembowski vill jag s�ga att r�det inte str�var efter en kompromiss .
. ( en ) fru talman ! jag vill f�rst tacka er alla f�r denna intressanta och v�rdefulla debatt .
�ndringsf�rslagen 1 , 6 , 7 och 8 g�ller ocks� v�gran till tilltr�de .
f�r att uppn� huvudsyftet med detta f�rslag , n�mligen att snabbt avveckla gamla oljetankfartyg med enkelskrov , �r vi beredda att g� med p� en strykning av det ekonomiska stimulanssystemet med differentierade hamn- och lotsavgifter .
medlemsstaterna m�ste f�rvissa sig om att det klassificeringss�llskap de v�ljer att arbeta p� deras v�gnar fullg�r uppgifterna till deras fulla bel�tenhet .
det l�mnar kvar �ndringsf�rslag 10 som g�ller den viktiga fr�gan om ansvarsbegr�nsningar .
jag vill avsluta med att p�minna om att f�r en m�nad sedan sj�nk ievoli-sun n�ra cherbourg med 6 000 ton farlig last .
" det �r naturligtvis t�nkbart att det n�gonstans sitter en inkompetent och provocerande tj�nsteman , men n�r femton l�nder godk�nner denna typ av svar , s� tycker jag , fru talman , att ni borde rikta en uppmaning till r�det att respektera det som �r en av parlamentsledam�ternas r�ttigheter .
bet�nkande ( a5-0342 / 2000 ) av ortuondo larrea fr�n utskottet f�r regionalpolitik , transport och turism om f�rslaget till europaparlamentets och r�dets direktiv om �ndring av r�dets direktiv 94 / 57 / eg om gemensamma regler och standarder f�r organisationer som utf�r inspektioner och ut�var tillsyn av fartyg och f�r sj�fartsadministrationernas verksamhet i f�rbindelse d�rmed ( kom ( 2000 ) 0142 - c5-0175 / 2000 - 2000 / 0066 ( cod ) )
om �ndringsf�rslag 2 :
( parlamentet antog resolutionen . )
skapandet av syssels�ttning m�ste f�rbli en av v�ra st�rsta prioriteringar .
samtidigt l�mnas de kapitalistiska rederiernas verksamhet okontrollerad genom att bekv�mlighetsflagg anv�nds och villkoren f�r den v�rldsomsp�nnande sj�farten f�rs�mras .
europeiska kommissionens f�rslag ser betryggande ut men �r inte tillr�ckligt skyddat mot v�lmedvetet motarbetande .
f�r att g�ra det m�ste vi f�rs�kra oss om att de �tg�rder vi i dag f�resl�r kommer att till�mpas av alla europeiska unionens medlemsstater .
kommissionen vill helt riktigt f�rebygga att europa hamnar p� efterk�lken gentemot amerika .
m�nga tekniker understryker i dag de sv�righeter man st�ter p� vid inspektion av utrymmet mellan de b�da skroven och underh�llet av detta utrymme .
det r�r sig om ett viktigt , men inte tillr�ckligt beslut .
dessutom har jag r�stat f�r alla de �ndringsf�rslag som f�rb�ttrar och sk�rper kommissionens f�rslag .
en �versyn av direktiv 94 / 57 / eg br�dskar , desto mer som malta och cypern �r ans�karl�nder , med v�rldens fj�rde respektive sj�tte st�rsta flotta .
det sparas in p� hamnavgifterna genom att segla vidare vid stormv�der och genom att �ven vid andra tillf�llen acceptera risken f�r att olyckor med d�dlig utg�ng kan intr�ffa .
sj�s�kerheten skall inte bara vara en fr�ga som tas upp i krissituationer , efter varje ny katastrof som drabbar v�ra kuster , utan omfattas av en integrerad och kontinuerlig politik p� internationell niv� .
lika lite bryr vi oss om ifall stadgan �ver grundl�ggande r�ttigheter inf�rlivas i eller h�lls utanf�r f�rdraget , f�r i alla h�ndelser v�grar denna stadga , som p�st�s g�lla grundl�ggande r�ttigheter , att ta upp arbetstagarnas element�ra r�ttigheter och �ppnar dessutom d�rren f�r socialt regressiva �tg�rder .
det ser jag som ett avg�rande kriterium f�r att bed�ma nicef�rdraget .
. ( fr ) inf�r toppm�tet i nice och utan att f�regripa resultaten av detta , vill jag ber�mma det franska ordf�randeskapets omfattande arbete och de flesta av ministrarna , som varken har sparat tid eller m�da f�r att regelbundet bes�ka v�rt parlament i utskotten och i kammaren .
debatten och den resolution europaparlamentet har antagit bidrar till allvarliga orosmoment om vad som skall beslutas under toppm�tet i nice , s�rskilt n�r det g�ller m�jliga sk�rpningar av restriktionerna f�r suver�niteten i sm� l�nder som portugal , f�r att st�rka federalismen och den milit�ra inriktningen p� f�rsvars- och s�kerhetspolitiken , och n�r det g�ller de svaga och klart otillr�ckliga �tg�rderna p� det sociala omr�det .
om f�rdragsreformen och utvidgningen skall bli framg�ngsrika m�ste de f� fullt st�d av folket .
de reformer som f�reslagits av parlamentsledamot malcolm harbour om vitboken �r reformer som styrs av sunt f�rnuft .
de v�ljare som jag h�r f�retr�der st�ller sig n�mligen inte bakom en enda av dess m�ls�ttningar .
det blir allt mer uppenbart att den p�b�rjade debatten om proportionaliteten ( vad avser r�ster i r�det och platser i europaparlamentet ) , det vill s�ga om maktf�rh�llandena mellan medlemsstaterna , har �ppnat en pandoras ask som det blir sv�rt att st�nga i nice .
s� om ni kan undvika krig , som ni har gjort hittills , s� skulle ni g�ra det viktigaste som n�gonsin har gjorts i hela v�rlden .
. ( fr ) delegationen f�r det andra europa inom gruppen unionen f�r nationernas europa har beslutsamt r�stat emot initiativbet�nkandet fr�n utskottet f�r utrikesfr�gor som f�rsvarades av brok .
jag har en systerson som har varit p� natos baser i usa f�r att l�ra sig flyga jaktplan , och han befordrades , han �r med andra ord redo att arbeta som pilot inom flygvapnet .
det �r upp till varje enskild medlemsstat att besluta om man vill delta i en gemensam europeisk s�kerhets- och f�rsvarspolitik .
vi �r �vertygade om att ett fredens europa inte skapas genom milit�rallianser .
vi beh�ver ingen euromilitarism .
. jag uppskattar f�rs�ket att utveckla en gemensam europeisk s�kerhetspolitik , men �r emot utvecklandet av ett gemensamt milit�rt f�rsvar .
vi anser inte att upprustning och d�rmed �kade milit�ra utgifter �r svaret p� europas utmaningar under denna era .
vi har 19 �verv�ganden och 23 punkter med 36 stycken .
men dokumentets spr�kliga form g�r ut�ver detta .
problem , som tas upp i bet�nkandet , kan l�sas med en human asyl- och flyktingpolitik , en arbetsorganisation som tar h�nsyn till balans mellan arbete och fritid samt genom ett solidariskt , samh�lleligt ansvarstagande f�r personer med s�rskilda behov .
f�redraganden anser att det kr�vs en r�ttslig ram p� europeisk niv� som g�r det m�jligt f�r personer som tillhandah�ller hush�llstj�nster att omfattas av en arbetarskyddslagstiftning .
hon vill att denna typ av arbete skall erk�nnas som ett yrke i sin egen r�tt och kr�ver att europeiska best�mmelser skall utarbetas om dessa arbetares r�ttigheter - f�r n�rvarande varierar situationen fr�n land till land .
bet�nkande ( a5-0327 / 2000 ) av guy-quint
sv�gerpolitik och bristande �ppenhet m�ste ocks� f�rsvinna inom kommissionens enheter , s�rskilt n�r det g�ller rekrytering av tillf�lligt anst�llda .
det �r d�rf�r l�mpligt att minuti�st vaka �ver att dessa �taganden respekteras i l�ngt st�rre utstr�ckning �n vad som tidigare skett .
jag r�stade f�r lamassoure-bet�nkandet som i f�rsta hand avser de institutionella aspekterna p� kommissionens reformering .
det beklagar jag och d�rf�r har vi ocks� som partigrupp avst�tt fr�n att r�sta , eftersom vi anser att det inte �r bra f�r de icke-statliga organisationerna .
fru talman ! f�r det andra skulle jag , med tanke p� den m�ngd motstridig information som vi har f�tt under dagens lopp , vilja att ni p� ett tydligare s�tt f�rklarar f�r kammaren hur strukturen p� diskussionen med det franska ordf�randeskapet avseende r�dets m�te i nice kommer att vara och p� vilket s�tt man kommer att presentera r�dets ordf�randes deltagande .
vill ni inte ha n�gon resolution ?
fru talman , ingen underskattar betydelsen och omfattningen av detta toppm�te som dessutom �r det l�ngsta toppm�tet i europeiska unionens historia .
konstitutionella fr�gor . ( it ) fru talman !
tack , herr h�nsch , f�r detta uppbyggliga bidrag .
fru talman ! mot bakgrund av det beslutet och eftersom kommission�r liikanen inte kommer att n�rvara p� torsdag men kan n�rvara p� onsdag , undrar jag om det skulle kunna vara n�jligt att tidigarel�gga fru gills bet�nkande om europeiskt digitalt inneh�ll fr�n torsdag till onsdag f�r att fylla den luckan .
fru talman ! i detta �gonblick , och sedan den 20 oktober , hungerstrejkar 200 politiska f�ngar till d�ds i turkiet f�r att protestera mot den politik som bedrivs av den turkiska regeringen vilken anv�nder de " vita " isoleringscellerna f�r att bryta ner f�ngarnas moral och motst�nd .
. ( nl ) fru talman ! det �r nu andra g�ngen i �r som vi diskuterar det h�r direktivet och �terigen har det l�mnats in m�nga �ndringsf�rslag .
trots denna tydliga linje m�ste vi inse att vi �r ett parlament i en union som hyllar r�ttsstatens principer och det inneb�r att vi m�ste erk�nna gr�nserna f�r v�r beh�righet , att vi m�ste veta hur l�ngt gr�nserna g�r f�r den beh�righet vi l�nar fr�n artikel 95 , den r�ttsliga grund vi �beropar f�r det nya tobaksdirektivet .
f�r att f�rsvara denna grundl�ggande princip f�reslog vi att den r�ttsliga grunden skulle ut�kas till att �ven omfatta artikel 133 i f�rdraget , men framf�r allt sk�t vi upp det datum f�re vilket medlemsstaterna m�ste till�mpa den till den 1 januari 2007 .
l�t oss vara absolut s�kra p� att de �r informerade n�r de fattar beslutet p� det ena eller andra s�ttet .
vi menar dock att det �r mycket stora skillnader mellan fr�gan om tobaksreklam och detta direktiv .
domstolen har n�mligen just upph�vt direktivet fr�n 1998 genom vilket reklam och sponsring av tobaksprodukter f�rbjuds .
r�dets f�rslag om texternas storlek p� andra f�rpackningar �n cigarettpaket tycker jag emellertid �r b�ttre �n det som st�r i �ndringsf�rslag 25 , eftersom gr�nsen 50 cm � ligger alldeles f�r n�ra hela ytan p� ett paket cigaretter .
detta �r det som bekymrar mig i denna fr�ga .
och d�rf�r har de en korrekt r�ttslig grund som utg�r fr�n tidigare artikel 100a eller den nuvarande artikel 95 .
dessutom �r jag r�dd f�r att det skall vara en d�lig f�rebild f�r att senare �ven s�tta varningstexter p� andra produkter .
herr talman ! det �r rimligt att s�ga att vi har en moralisk skyldighet att fullt informera de 30 miljoner konsumenterna i europeiska unionen om cigaretters risker f�r folkh�lsan .
s� i st�llet f�r att exportera cigaretter kommer vi att exportera jobb - 4 000 av dem i min region enbart .
herr talman ! jag vill f�rst och fr�mst gratulera maaten till ett lysande bet�nkande .
herr talman ! r�kning �r v�r tids tragedi - den st�rsta orsaken till sjukdomar som kan f�rebyggas i hela europeiska unionen .
om ni anf�r artikel 133 f�r exportf�rbudet , kan ni konstatera att det inte �r en uppgift f�r en gemensam handelspolitik att diktera ett tredje land vad man sj�lv skall importera .
det f�r inte bli n�got undantag f�r m�rkning annars kommer vi bara att skapa nya missf�rh�llanden inom konkurrens och den inre marknaden .
jag hoppas att kommission�ren kan utlova en f�rst�rkning av personalst�det inom kommissionen .
herr bowis fr�gade om undantaget skulle g�lla .
de fastslog vidare i punkt 117 i domen : " det har ovan i punkterna 98 och 111 i denna dom p�pekats att artikel 100a i f�rdraget skulle kunna m�jligg�ra antagandet av ett direktiv som f�rbjuder vissa former av reklam f�r och sponsring till f�rm�n f�r tobaksvaror .
kommissionen skulle f�redra att granska den tillg�ngliga informationen och rapportera tillbaka i vederb�rlig ordning .
kommissionens rapporter om till�mpning av punktskattedirektiven hanterar detta problem p� l�mpligt s�tt .
som f�redragande skulle jag rekommendera att dessa �ndringsf�rslag st�ds d� de verkar mycket f�rnuftiga .
den timme av extra dagsljus som erh�lls genom �verg�ngen till sommartid gynnar i synnerhet sektorerna f�r turism och fritidsaktiviteter som har f�tt f�rnyad verksamhet i direkt samband med de ljusare och l�ngre kv�llarna .
jag har sagt det f�r att min fraktion och �ven jag �r �vertygade om att europa har st�rre problem och uppgifter .
de �ndringsf�rslag som v�ckts av parlamentet och f�redraganden �r d�rf�r - enligt min �sikt - inte till hj�lp eftersom de snarare medf�r os�kerhet �n �kat f�rtroende .
till exempel f�r transportsektorn i synnerhet men ocks� andra industrisektorer , beh�ver en stabil , l�ngsiktig planering beroende p� tekniska krav i samband med planl�ggning av tidsscheman f�r transporter .
n�sta punkt p� f�redragningslistan �r andrabehandlingsrekommendationen ( a5-0349 / 00 ) av liese f�r utskottet f�r milj� , folkh�lsa och konsumentfr�gor om r�dets gemensamma st�ndpunkt inf�r antagandet av europaparlamentets och r�dets direktiv om tilln�rmning av medlemsstaternas lagar och andra f�rfattningar r�rande till�mpning av god klinisk sed vid kliniska pr�vningar av humanl�kemedel ( 8878 / 1 / 2000 - c5-0424 / 2000 - 1997 / 0197 ( cod ) ) .
n�r det g�ller den direkta nyttan , m�ste man vid kliniska f�rs�k skilja mellan medicinering och �tf�ljande unders�kningar , som �r n�dv�ndiga f�r att dra slutsatser f�r kommande patienter .
of�rm�gna vuxna f�r avslutningsvis bara delta i de pr�vningar som avser den sjukdom som de lider av och �r ursprung till deras of�rm�ga .
n�gra ord om en annan mycket viktig fr�ga i mina �gon , jag vill tala om �ndringsf�rslag 30 som r�r icke kommersiella kliniska pr�vningar .
av den anledningen b�r l�karvetenskapen ha alla medel att tillg� f�r en h�g grad av skydd f�r den personliga h�lsan och f�r folkh�lsan .
jag f�rklarar debatten avslutad .
vi b�r inte gl�mma att gemenskapens regelverk som g�ller dessa program i sj�lva verket kommer att �verf�ras till det nya h�lsoprogrammet vilket utarbetas f�r n�rvarande , s�ledes �r det r�tt att de f�rl�ngs .
jag tror inte , s�som trakatellis sade , att man kan leka med de sjuka personers h�lsa , som v�ntar p� v�r hj�lp , och med de icke-statliga organisationer som beh�ver dessa gemenskapsanslag f�r att sk�ta folkh�lsopolitiken ute p� f�ltet .
programmen f�r att f�rhindra narkotikaberoende m�ste ocks� inriktas inte bara p� krisomr�den utan p� m�nga andra omr�den inom europeiska unionen .
sammanfattningsvis , fru talman , m�ste jag s�ga att utvecklingen inom folkh�lsosektorn i europeiska unionen g�r f�r l�ngt f�r mig .
brottsoffrets st�llning i det straffr�ttsliga f�rfarandet
jag vill ocks� understryka att trots dess betydelse och att den �r en obligatorisk referenspunkt i europa s� har konventionen �nnu inte ratificerats ( den 18 september 2000 ) av f�ljande medlemsstater i europeiska unionen : �sterrike , belgien , grekland , irland , italien , portugal och spanien .
den andra aspekt som spelat en viss roll , var fr�gan om videof�rh�r .
vi har kanske �gnat f�r lite tid �t brottsoffren , vilka oftast �r den svagaste delen i denna v�rld .
slutligen �r detta beslut viktigt eftersom parlamentet har m�jlighet att f�rb�ttra lagf�rslaget betydligt genom just cerdeiras utm�rkta bet�nkande , som utskottet f�r medborgerliga fri- och r�ttigheter har inst�mt i .
dessutom konstateras det att brottsoffer bem�ts diskriminerande vid anm�lan av brott .
den skyldige , arturo lojacono , har identifierats och d�mts , men flydde utomlands .
det kan vara sv�rt f�r ett utl�ndskt brottsoffer att p� avst�nd f�lja de r�ttsliga f�rfarandena , och det �r klart att det d� beh�vs s�rskilda �tg�rder .
den var f�rem�l f�r sv�ra diskussioner i r�det .
kommissionen �nskar forts�tta unders�kningen av genomf�rbarheten av ett s�dant projekt .
herr posselt , vi kommer att vidarebefordra era synpunkter till kvestorskollegiet f�r att de skall fatta det beslut som de anser vara l�mpligast och att detta kommer till samtliga ledam�ters k�nnedom .
kommissionen st�der d�rf�r r�dets anh�llan om br�dskande f�rfarande och ber europaparlamentets ledam�ter v�nligast om st�d f�r detta br�dskande f�rfarande .
jag har h�rt av min ordf�rande i budgetutskottet att det faktiskt skulle vara f�rsta g�ngen som ett enande uppn�tts mellan r�det och parlamentet i en f�rlikning .
kommissionen har lagt fram sin rapport med analysen av de utest�ende �tagandena och deras strategiska ansats f�r att uppl�sa les restes � liquider .
vi kan finansiera samarbetet med den baltiska regionen och v�ra krishanteringsstyrkor , och vi har utrustat meda med 40 miljoner euro mer �n r�det hade avsett .
eftersom jag bara f�tt s� lite tid till f�rfogande , vilket jag beklagar s�tillvida som budgeten �ven f�r f�redragandena hade f�rtj�nat mer �n de skrattretande tv� och en halv minuterna , m�ste jag inskr�nka mig till n�gra f� p�pekanden .
. ( es ) herr talman ! n�r en delegation fr�n detta parlament bes�kte folkrepubliken kina f�r en tid sedan var vi i xiamen i den syd�stra delen av landet , och vi s�g d�r en � i horisonten .
de tre institutionernas f�retr�dare sparade inte p� anstr�ngningarna n�r det g�llde att uppn� en total �verenskommelse om budget 2001 och jag vill i detta sammanhang framf�ra r�dets tack s�v�l till ledam�terna i den parlamentariska delegationen som till fru schreyer .
det gl�der mig att v�ra institutioner lyckats komma �verens om att vid en enda behandling anta samtliga best�ndsdelar i denna �ndringsskrivelse nr 2 som inte bara g�ller jordbruksutgifterna utan �ven fiskeriavtalen och inf�randet av ett prelimin�rt saldo f�r budget�ret 2000 i den ursprungliga budgeten f�r 2001 .
jag f�ster f�r min del mycket stor betydelse vid den .
efter denna �versikt vill �ven jag betona det utm�rkta klimat i vilket detta budgetf�rfarande genomf�rts .
det �r ur kommissionens synpunkt det faktum att den andra pelaren i jordbrukspolitiken , n�mligen st�det till landsbygdens utveckling , uppvisar den st�rsta �kningen . h�r uppg�r �kningen till 10 procent , och det anser jag v�rt att p�peka , ty d� st�r totalt sett 4,5 miljarder euro till f�rfogande .
. ( fr ) herr talman ! jag skulle vilja svara colom i naval p� fr�gan om utnyttjandet av mekanismen f�r flexibilitet n�r det g�ller �versynen av budgetplanen .
vi ber�mde kommission�r busquin , som har �vertr�ffat v�ra f�rv�ntningar p� det omr�det .
herr talman ! som f�redragande av yttrandet fr�n utskottet f�r utveckling och samarbete vill jag f�r det f�rsta konstatera att europaparlamentet vunnit en stor seger genom att inbesparingen p� latinamerikanska , asiatiska och afrikanska fattigdomsprogram har upph�vts .
i synnerhet vill jag n�mna euronews s� att m�nniskor kan se i pressen vad parlamentet och unionen arbetar med .
vi har en budget som �r under 1,06 procent , vi har en budget , herr colom , som ligger inom ramen f�r budgetplanen .
jag vill tacka fru schreyer , som ocks� har hj�lpt oss vidare med sitt mycket konstruktiva s�tt att ta itu med saker och ting , och naturligtvis ocks� min v�n jutta haug , som har �stadkommit ett utm�rkt arbete , och likas� joan colom i naval och �ven markus ferber .
ni s�ger hela tiden att budgetplanen �r okr�nkbar f�r er .
�ven v�r grupp kommer att r�sta f�r denna budget , eftersom den visar att vi trots �kande problem p� ett f�red�mligt s�tt �ter har skapat en kompromiss .
k�ra kolleger ! vi v�lkomnar nu jacques chirac , republiken frankrikes president och unionens tj�nstg�rande ordf�rande ,
man m�ste ocks� v�lkomna den europeiska andan som slutligen gjorde det m�jligt att l�mna nice efter att ha l�st de fr�gor som f�rblev ol�sta i amsterdam och efter att ha f�rberett framtiden .
jag kommer nu till ett av de mest positiva resultaten av regeringskonferensen .
f�r utvidgningen �r verkligen europas stora fr�ga .
man kommer i framtiden att bed�ma hela dess omfattning och jag hyllar er kammare som i h�g grad bidragit till att den kunnat utarbetas .
f�r ett �r sedan sj�nk erika utanf�r frankrikes kust . trots den fantastiska insatsen fr�n frivilliga och de offentliga myndigheterna lider kusten fortfarande av konsekvenserna av f�rlisningen .
till att b�rja med avslutade vi i nice den cykel som inleddes vid europeiska r�det i k�ln och helsingfors .
man kan gl�djas �t att unionen kunnat avisera att den skulle avs�tta cirka 13 miljarder euro under sju �r , inbegripet naturligtvis l�nen fr�n europeiska investeringsbanken .
n�r det g�ller utvidgningen , s� har den strategi som kommissionen f�reslog godk�nts . dessutom godk�nde r�det den sociala dagordningen , resultatet av ett fruktbart samarbete med ordf�randeskapet , vilket redan har p�pekats h�r .
parlamentet uppn�r framf�r allt att det bildas europeiska politiska partier . kommissionen f�rsvarade - dessv�rre utan framg�ng , men debatten �r inte avslutad - v�r gemensamma str�van att skydda unionens ekonomiska intressen genom f�rslaget att tills�tta en allm�n �klagare .
vi har tyv�rr under de senaste m�naderna - och inte heller detta f�r n�gonsin upprepas , eftersom det verkar som ett smygande gift i europeiska unionen - upplevt motsatsst�llningen mellan de stora och de sm� l�nderna , varvid flera stora l�nder har upptr�tt mycket sm�aktigt , och flera sm� l�nder har upptr�tt storartat .
det handlar om en tillbakag�ng som kommer att f� �terverkningar inom alla omr�den inom gemenskapen och jag f�rutsp�r , herr ordf�rande f�r europeiska r�det , att v�ra medborgare - och �ven parlamentarikerna och regeringscheferna �r jag r�dd - kommer att bli tvungna att s�tta sig i skolb�nken igen f�r att f� undervisning om matematiska kalkyler .
jag kan s�ga att det finns delar som vi tycker bra om och mycket som ber�r oss .
( appl�der )
det stora antalet blockeringar mellan de femton medlemsl�nderna under toppm�tet �r symptomatiska .
utan folkligt st�d , eftersom det inte finns n�got europeiskt folk , tvingas staterna av sin allm�nna opinion att p� ett allt mer envist s�tt f�rsvara sina nationella intressen , med risk f�r att �ndra det maximala antalet ledam�ter i europaparlamentet som fastst�llts i amsterdamf�rdraget som redan �r f�r�ldrat , med risk f�r att �ka antalet kommission�rer till 27 , trots att den nuvarande kommissionen med femton ledam�ter inte fungerar .
i vilken situation kommer alla dessa m�nniskor att ha dragit in frankrike , n�r den europeiska bubblan spricker och fransm�nnen bara har den bittra smaken kvar i munnen av att �nnu en g�ng ha l�tit sig luras av medelm�ttiga och intresserade ledare ?
bakom detta finns snarare graverande problem och oro och alltid resultatet av nationell opinionsbildning , som man inte f�r skjuta �t sidan , utan m�ste ta p� allvar .
ordf�randeskapet har beklagat denna otillr�cklighet . ordf�randeskapet hade sj�lvt f�rbeh�ll och kr�vde en stor anstr�ngning f�r att frankrike skulle g�ra framsteg inom omr�den som var s�rskilt k�nsliga f�r landet .
d�rf�r f�religger dessa �ndringsf�rslag , de s� kallade kompromiss�ndringsf�rslagen , fr�n tre grupper .
det var n�dv�ndigt att finna en l�sning p� m�ngfalden juridiska och administrativa situationer som till�mpas p� kliniska f�rs�k i medlemsstaterna .
jag tror att det skulle vara r�tt att ocks� och slutgiltigt f� en sommartid som �r densamma i samtliga stater i europeiska unionen . "
nu kommer vi till r�stf�rklaringarna om cerdeira mortereros bet�nkande .
l�mpliga �tg�rder m�ste vidtas f�r att ge brottsoffer f�ljande r�ttigheter : att tillhandah�lla och f� information ; kommunikationsm�jligheter ; deltaga i f�rfarandet och tillg�ng till gratis r�ttshj�lp ; en l�mplig niv� av skydd och privatliv ; m�jlighet att ans�ka om ers�ttning inom brottsm�lf�rfarandet och att f� en tvist bilagd genom f�rlikning .
europeiska r�det / franska ordf�randeskapet ( forts�ttning )
det f�rklarar varf�r m�nga av oss tyckte att nice var helt hoppl�st .
stats- och regeringscheferna har just erk�nt i nice det vi sade efter amsterdam , att metoden med regeringskonferensen inte l�ngre lyckas utveckla europa p� ett positivt s�tt .
som f�retr�dare f�r de partier som f�renats i europeiska fria alliansen vill jag varna fr�mst r�det men �ven kommissionen f�r om eu inte vill vara mer �n ett mellanstatligt f�rbund .
herr talman ! det n�gorlunda samst�mmiga budskapet fr�n r�dsordf�randen , kommissionen och regeringscheferna g�r ut p� att nicef�rdraget garanterar ramarna f�r ett samlat europa .
det inneb�r att det demokratiska underskottet �ter har blivit st�rre .
l�t oss se seri�st p� det som har h�nt .
i sj�lva verket �r det presidenten som �r orealistisk , om han tror att det med ett s�dant f�rdrag skall bli m�jligt att utvidga unionen .
herr talman ! m�tet i nice var och borde vara ett historiskt m�te , ett startskott f�r det nya europa , det nya seklets europa , det stora europa , ett europa f�r alla europ�er .
utvidgningen har st�llt er och oss alla inf�r samma uppgift som monnet och schuman och andra f�r femtio �r sedan stod inf�r : n�mligen att utveckla en metod , en struktur och en vision f�r europas framtid .
�terst�r s�ledes bara ett litet gl�dje�mne : utvidgningen .
det framtr�der fyra huvudproblem .
denna passus ansluter sig till europaparlamentets uppfattning att europeiska unionen inte kan utvecklas vidare genom den hittillsvarande metoden med regeringskonferenser .
ocks� jag f�rs�ker - liksom frankrikes president h�r i f�rmiddags - t�nka mig vad som skulle ha h�nt om vi hade kommit hit utan nicef�rdrag .
vi f�rs�kte arbeta p� en princip med enkel r�stviktning , inom denna om�jlighet , och jag tror att resultatet totalt sett �r r�ttvist .
vi f�r sedan alla tillsammans se hur vi skall g�ra f�r att forts�tta .
vi m�ste avskaffa regeln med konsensus , �ven i ett framtida konvent .
i samtliga dessa fall drog vi slutsatsen att dessa f�rdrag inte var helt tillfredsst�llande , inte svarade mot alla v�ra f�rhoppningar men trots det utgjorde ett steg fram�t och �tminstone var b�ttre �n status quo .
m�nga m�nniskor som granskar f�rdraget fr�n nice kommer att undra varf�r det utformades p� det s�ttet .
men europeiska r�det i nice inneb�r , som s� m�nga andra toppm�ten i europeiska unionens historia , en triumf f�r verkligheten och en triumf f�r pragmatismen �ver utopin .
vi skulle med b�ttre samvete ocks� ha kunnat f�rmedla ett b�ttre och starkare europeiskt resultat till befolkningen .
detta toppm�te skulle ha varit en fullst�ndig framg�ng om den n�dv�ndiga �versynen av f�rdragen kr�nts av samma succ� som de kapitel jag just n�mnt .
dessutom �r det mer demokratiskt .
blair �terv�nde till storbritannien som en vinnande hj�lte f�r att han inte hade avst�tt det h�r , inte hade avst�tt det d�r och hade k�mpat f�r storbritanniens intressen .
i dagens debatt har vi inte dolt tillfredsst�llelsen �ver och , i �nnu h�gre grad , missn�jet med nicef�rdraget , ibland av olika sk�l men med samma k�nslor och med samma oro .
en bra signal till v�ra partner i s�der .
det st�mmer att v�r kammare snarare �r glest befolkad . men budgetdebatten har tyv�rr tagit l�ngre tid �n planerat och vi f�r inte , vare sig jag sj�lv eller de talare som f�ljer efter mig , m�jlighet att ta upp fr�gan med ordf�randeskapet .
herr talman , mina damer och herrar ! n�r budgeten st�lldes upp tog man h�nsyn till principerna sparsamhet , social och ekonomisk balans .
l�t oss inte lura oss sj�lva , detta �r en bra budget .
det som vi talar om �r ett system f�r f�rtidspensionering , vilket �nnu inte har n�gon r�ttslig grund ; ingen vet om det som kommer att f�resl�s skall vara obligatoriskt eller ej obligatoriskt och det �r trots allt ett p.m. som st�r p� spel .
herr talman , mina damer och herrar , fru kommission�ren , r�dets f�retr�dare , mina damer och herrar , �rade f�redragande ! under varje budget�r vinner parlamentet budgetf�rdelar .
och jag g�r lite l�ngre , f�r det r�cker n�mligen inte med att bara ha kr�vande och genomblickbara regler vid verkst�llandet av budgeten , som annulleringen av �taganden efter tv� �r av l�g genomf�randegrad .
det k�nner vi alla till .
det �r lagrar som vi delar ut i f�rskott , och ni kan vara s�kra p� att vi i framtiden kommer att f�rs�ka kontrollera det str�ngt .
h�r har ni nu ocks� �tg�rder som uttryckligen fr�mjar milj�skyddet .
. ( nl ) herr talman ! f�rbindelserna med ryssland har �ndrats i grunden sedan det kalla krigets dagar .
jag anser f�r �vrigt att rysslands intressen inte m�rks riktigt i budgeten , men i det avseendet tycker vi annorlunda �n socialdemokraterna .
nu �r jag positiv till att uppmuntra ryssland och ukraina att g� i v�r riktning och samarbeta med andra alliansl�nder i krishanteringsinsatser , men jag skulle inte vilja att vi g�r i deras riktning eller att vi anpassar v�r politik f�r att foga oss efter dem .
om denna situation inte snarast �ndras genom att man i ryssland skapar den n�dv�ndiga r�ttsliga och s�kerhetsm�ssiga ramen och p� s� vis �stadkommer ett v�nligare investeringsklimat , d� finns det trots de nya h�ga priserna p� mineralolja knappast n�gon utv�g ur den ekonomiska krissituationen .
det betyder att vi har ett gemensamt ansvar f�r freden i kaukasus , f�r milj�skyddet i ryssland och f�r den inhemska befolkningen d�r .
jag anser att l�sningen inte kan vara milit�r , att situationen visar det tillr�ckligt och att l�sningen bara kan vara politisk .
nyligen hamnade den k�nda ryska oppositionspolitikern grigorij jawlinskij i de v�sterl�ndska tidningarna igen .
kreativa l�sningar f�r befolkningen i kaliningradomr�det , med tanke p� deras kommande frihet till transitresor genom litauen och polen , b�r ocks� f�rdigf�rhandlas f�re polens och litauens anslutning till eu .
det �r inte bara f�r att alla europeiska stormakter framf�r allt vill f�rsvara intressena hos sina egna kapitalistiska grupper , men vad har egentligen det kapitalistiska europa att erbjuda ryssland ?
den dubbelstrategi som oostlander f�resl�r , och som f�rtj�nar ber�m , erbjuder en utv�g .
hans bet�nkande har v�lkomnats av alla delar av parlamentet utom kanske av dem som ser tillbaka med nostalgi till de inte s� gyllene tiderna som bevaras i minnet av ett stort antal modiga , sovjetiska avhoppare .
jag �r angel�gen att f� arbeta i n�ra samarbete med det tilltr�dande svenska ordf�randelandet f�r att skapa konkreta framsteg med den nordliga dimension .
det �r p� grund av att vi anser v�rt f�rh�llande med ryssland s� viktigt som dessa fr�gor �r viktiga .
ang�ende : genetiskt modifierade organismer och gr�dor sedan v�ren 2000 har man i olika l�nder i eu kunnat konstatera flera fall av genetiskt modifierade organismer och gr�dor - bomull , raps och majs - som sl�ppts ut i milj�n .
i denna gemensamma st�ndpunkt �l�ggs medlemsstaterna mycket str�ngare skyldigheter .
det skulle fr�n r�dets sida vara b�de of�rsiktigt och dumt .
f�r det andra : har r�det l�tit sig informeras av europar�dets kommissarie med ansvar f�r de m�nskliga r�ttigheterna , som ju �r v�l f�retr�dd p� ort och st�lle ?
r�dets ordf�rande m�ste �nd� veta om han har tr�ffat masjadov eller inte .
vilka �ndringar har r�det f�r avsikt att tillf�ra direktivet i fr�ga ( 92 / 12 / eeg ) s� att ansvaret mellan avs�ndare och mottagare kan delas upp med precision och m�jligheterna till bedr�geri undanr�jas ?
denna rapport visar , som ni s� riktigt s�ger , att skattebedr�geriet i gemenskapen n�tt en oroande niv� .
jag skulle vilja f�sta den �rade parlamentsledamotens uppm�rksamhet p� det faktum att det i f�rslaget till direktiv faktiskt n�mns , i sk�l 3 , att dess till�mpning inte p�verkar �taganden enligt gen�vekonventionen av den 28 juli 1951 om flyktingars status , s�som den �ndrats genom new york-protokollet av den 31 januari 1967 .
. ( fr ) det f�rslag till r�dets f�rordning som kommissionen nyligen lagt fram om �ndring av r�dets f�rordning ( eg ) nr 2820 / 98 f�r att utvidga tullfriheten till produkter fr�n de minst utvecklade l�nderna utan n�gon kvantitativ begr�nsning kommer av gemenskapens initiativ som syftar till att f�rb�ttra de minst utvecklade l�ndernas tilltr�de till marknaden .
. ( fr ) jag skulle bara vilja f� er att f�rst� , eftersom det �r mitt sista m�te h�r , vad det h�r momentet best�r i .
avslutningsvis kan icke testade djur som �r �ldre �n trettio m�nader inte l�ngre ing� i livsmedelskedjan .
som ni sj�lv betonade �r det dj�rva beslut , som nyligen fattats eftersom det senaste jag n�mnde �r fr�n den 4 december , allts� f�r en vecka sedan .
partiet �nskar f�rena islam och modernitet och skulle i h�g grad kunna bidra till att ge ny fart �t den demokratiska utvecklingen , vilken minst sagt avstannat , och f�ljaktligen till att konsolidera r�ttsstaten . ett f�rbud har utf�rdats mot detta parti med den f�rlegade f�rev�ndningen att det utg�r ett hot mot statens s�kerhet .
ang�ende : fn : s specialsession om barn fn : s generalf�rsamlings specialsession om barn i september 2001 kommer att diskutera barnens situation i v�rlden och man har f�r avsikt att anta en ny handlingsplan f�r att se till att barnens r�ttigheter f�rverkligas i hela v�rlden .
fr�ga nr 11 fr�n ( h-0894 / 00 ) :
loizidou-fallet : tv� f�llande domar mot turkiet .
detta sker framf�rallt i f�ngelset longuenesse i frankrike och g�ller l�ngtradarchauff�rer fr�n f�renade kungariket och andra l�nder .
i enlighet med artikel 23 i f�rdraget om europeiska unionen antar r�det detta beslut enh�lligt , vilket f�r �vrigt g�ller samtliga �vriga beslut som f�r konsekvenser f�r f�rsvarsomr�det .
fr�ga nr 22 fr�n ( h-0918 / 00 ) :
som ni vet noterades tyv�rr inga framsteg i nice p� detta omr�de .
herr talman , efter f�r�ndringarna och den demokratiska utvecklingen i jugoslavien , stabiliserings- och associeringsavtalet mellan europeiska unionen och f.d. jugoslaviska republiken makedonien och efter det f�rest�ende stabiliserings- och associeringsavtalet med republiken kroatien ser det ljust ut f�r demokratiseringen och normaliseringen p� v�stra balkanhalv�n , och i synnerhet kroatien kan spela en avg�rande roll i denna riktning .
�ven den �ndrade attityden fr�n de nyvalda kroatiska myndigheternas sida till internationella krigsf�rbrytartribunalen f�r f.d. jugoslavien r�knas kroatien till godo .
jag vill ocks� betona att kroatien bem�dar sig att f� fullst�ndig ordning p� sina f�rbindelser med grannl�nderna .
detta land hade till skillnad fr�n grannlandet slovenien inte omedelbart efter oberoendet �r 1991 kunnat utvecklas s� att det redan nu �r ett kandidatland .
. ( en ) herr talman ! jag �r glad att f� ge synpunkter p� det utm�rkta bet�nkandet av den �rade ledamoten baltas - framtagen , som flera �rade ledam�ter har sagt , med avsev�rd skyndsamhet - om kommissionens genomf�rbarhetsstudie om ett stabiliserings- och associeringsavtal med kroatien .
i f�rra m�naden , som kammaren k�nner till , var kroatien med ytterst imponerande effektivitet och diplomatisk fink�nslighet v�rd f�r det historiska toppm�tet i zagreb .
vi v�lkomnar parlamentets st�d hittills , inte minst f�r den viktiga fr�gan om r�ttslig grund f�r stabiliserings- och associeringsavtalen .
v�gen till demokrati , till respekt f�r m�nniskans r�ttigheter , till en bra regim- och r�ttsprincip , till utrotandet av korruptionen , verkar vara en l�ng v�g med m�nga hinder .
f�rra veckan togs 100 studenter till f�nga och fyra av dem l�mnades d�da tillbaks till deras f�r�ldrar .
eu-ambassaden i jakarta kan p�ta sig den samordningen .
( pt ) herr talman ! den positiva utveckling vi har sett i indonesien �r odiskutabel och detta g�r det tillr�dligt att skapa nya f�rbindelser och ett effektivt samarbete med detta land .
mer �n 100 000 flyktingar finns i v�stra timor och dessa anv�nds som m�nskliga sk�ldar av de moraliska och materiella anstiftarna till brotten i �sttimor .
p� m�nga platser �vertr�ffar v�ldet dialogen .
den internationella gemenskapen m�ste st�lla jakarta under maximal press f�r att f� slut p� v�ldet p� moluckerna .
jag anser att indonesien �r ett betydelsefullt land , men det st�r inf�r ett v�gval och det beror p� det internationella samfundets och europeiska unionens anstr�ngningar att i detta v�gval peka mot demokratin , mot respekten f�r de m�nskliga r�ttigheterna och mot r�ttsstaten , i annat fall kommer oordningen att f�rv�rras .
den st�ndpunkt vi m�ste ha r�rande indonesiens territoriella integritet �r enkel : vi m�ste f�lja internationell lagstiftning och f�renta nationernas resolution 2504 fr�n december 1969 .
herr talman ! jag v�lkomnar detta bet�nkande , men det k�nns en smula optimistiskt .
ett s�rskilt fall �r fortfarande den ol�sta fr�gan om v�sttimor .
det st�d som vi f�r n�rvarande ger justitieministern i jakarta �r avsett att hj�lpa honom i hans f�rs�k att bek�mpa korruption .
utvidgningen av gemenskapen och inf�randet av euromynten kan medf�ra ytterligare risker .
jag tackar kommissionen f�r dess anstr�ngningar och insatser ...
jag �r s�ker p� , fru kommission�r , att om man tar detta f�rsta steg , s� f�rlorar diskussionen om den europeiska �klagarmyndigheten karakt�ren av ett religionskrig mellan motst�ndare och f�respr�kare , vilket hittills har hindrat alla framsteg .
�ven om vi har all t�nkbar sympati f�r f�redraganden , fru theato , och hennes duktiga insatser f�r �vrigt , mots�tter vi oss inr�ttandet av en oberoende europeisk �klagarmyndighet , d�rf�r att den �r ett led i det federala europa som vi �r motst�ndare till .
herr talman ! det �r alltid ett n�je att tala efter dell ' alba f�r han f�r en brittisk euroskeptiker att l�ta mycket klok p� denna plats .
jag vill gratulera fru theato f�r hennes bet�nkande och i synnerhet f�r att hon anstr�ngt sig att komma hit , eftersom jag vet att hon inte k�nner sig s� bra i kv�ll .
strategin omfattar fyra handlingsomr�den : lagstiftningen betr�ffande bedr�geribek�mpning , det operativa samarbetet mellan de ansvariga myndigheterna , de interinstitutionella tillv�gag�ngss�tten f�r att bek�mpa bedr�gerier i tj�nsten och vidareutvecklingen av den straffr�ttsliga dimensionen .
n�sta m�l �r �r 2004 , n�sta regeringskonferens .
detta har h�nt vid flera tillf�llen avseende strukturfonderna exempelvis .
det �r ocks� ytterst viktigt att vi h�ller fast vid det ansvarsomr�de som kr�vs av oss och att vi i v�rt ansvarsfrihetsf�rfarande inriktar oss uteslutande p� det aktuella �ret .
n�gon g�ng m�ste vi �ndra p� r�dets st�ndiga fr�nvaro och dess oskyldiga attityd , r�det som aldrig b�r skulden f�r n�gonting .
revisionsr�tten redovisar rapporter och en av de viktigaste kunderna f�r de rapporterna �r parlamentet .
andemeningen i bet�nkandet �r , okonventionellt uttryckt , att budgetkontrollutskottet i framtiden kommer att kontrollera noggrannare och �ven vill ha noggrant besked om vart de europeiska skattepengarna har tagit v�gen .
jag fick h�ra - och det �r inte en isolerad h�ndelse - att i f�renade kungariket sade socialministern p� tv att om han kunde stoppa bedr�geriet skulle han kunna spara 6 miljarder gbp .
efter h�ndelserna f�rra �ret �r ert m�l att budgetkontroll- och ansvarsfrihetsf�rfarandet skall bli �ppnare och framf�r allt mer effektivt .
�ven detta m�ste man d� ta h�nsyn till .
den gemensamma st�ndpunkt som f�religger och som vi i dag skall besluta om anser jag har en hel rad avg�rande brister , som f�r �vrigt under debatten hittills principiellt sett inte har bestridits av n�gon .
om man reglerar n�got s�dant fr�n tre h�ll , d� �r det klart att det finns tillr�ckligt m�nga h�llpunkter och anledningar till tvister och att man d�rigenom inte skapar n�gon r�ttss�kerhet .
den europeiska enhetliga marknaden �r en paneuropeisk marknadsplats , men d�r b�rsmarknaden m�ste behandlas likadant som andra marknader s� att nationella gr�nser , �ven om de markerar olika r�ttsliga beh�righetsomr�den , inte inkr�ktar p� den �verensst�mmelse mellan regler som kr�vs p� hela marknadsplatsen .
det andra blocket innefattar en rad �ndringsf�rslag som syftar till att f�rb�ttra de anst�lldas delaktighet vid ett offentligt uppk�pserbjudande .
i f�rslagen finns tre viktiga element i ett skede d� det sker en f�r�ndring av vem som kontrollerar ett f�retag : skydd av minoritetsaktie�gare , �ppenhet om information r�rande ett uppk�pserbjudande och reglerande �vervakning av processen .
detta �r en fr�ga d�r tydlighet �r ytterst viktig .
man m�ste visa st�rre f�rst�else f�r de nationella s�rdragen , annars kan det f� f�r�dande konsekvenser f�r ett enskilt medlemslands f�retagsstruktur .
bolkestein har sj�lv sagt att det �r mycket viktigt att ledningen f�r uppk�pshotade f�retag samr�der med aktie�gare i detta fall .
herr talman ! det �r intressant att lyssna p� herr martin som engelsk talare och jag kan f�rs�kra honom att saker h�ller verkligen inte p� att rasa samman i den brittiska ekonomin �ven om mitt parti skulle se en ny regering .
det �ndringsf�rslaget syftar till att inf�ra ett instrument som g�r det m�jligt f�r en majoritetsaktie�gare att �verta �vriga v�rdepapper .
vi kan i det avseendet l�ra oss mycket av situationen i f�renta staterna och det borde mana oss till st�rre f�rsiktighet .
jag �r skyldig kollegerna dehousse och echerer stort tack , som i m�nga samtal har bidragit till de b�rkraftiga kompromisserna .
de bet�nkligheter som framf�rts fr�n olika h�ll kan sammanfattas i tv� stora grupper .
herr talman ! f�r att besvara det lyckade uttrycket fr�n den europeiska sammanslutningen av f�rfattar- och komposit�rsf�reningar , har det f�rslag vi diskuterar under granskningen i r�det varit f�rem�l f�r orimliga angrepp .
jag kommer att i mitt land tvingas arbeta h�rt f�r att �vertyga dem , men jag �r fast �vertygad om att harmoniseringen av f�ljer�tten , som europaparlamentet ser den , medf�r f�rdelar f�r alla ber�rda parter .
det har ingenting att g�ra med nationella s�rintressen , utan det har att g�ra med att bidra till en �ppen politisk diskussion .
med en artikel skulle det ha varit v�ldigt sv�rt att hitta konstn�rens familj ; enbart efterforskningsbyr�er och inkasseringsfirmor skulle ha dragit n�gon nytta .
den andra viktiga fr�gan �r taket som avskaffas i ert �ndringsf�rslag 7 .
jag noterar det .
denna viktiga fr�ga - som �r central f�r utskottet - b�r enligt min mening debatteras i dag .
det som har �verraskat mig n�got som f�redraganden i de senaste m�nadernas debatt �r att vi har f�rlorat dessa tre saker ur sikte .
utan att ifr�gas�tta moderniseringen och konkurrensuts�ttandet av alla postf�retag , m�ste medlemsstaterna forts�tta att skydda sina n�tverk av postkontor med personlig betj�ning i landsbygdsomr�den , en faktor som minskar avst�nden fr�n de perifera omr�dena till beslutscentrumen och d�rmed �r n�dv�ndig f�r den sociala sammanh�llningen av de minsta samh�llena och landsbygden .
det finns ingen anledning till att den tj�nst som erbjuds folken inte skall omfatta alla tekniska och ekonomiska framsteg . det faktum att man avskaffar speciella tj�nster tror jag d�rf�r �r ett framsteg mer �n ett klarg�rande .
�rade fru talman , �rade herr kommission�r ! jag vill b�rja med att tacka v�r kollega markus ferber � min grupps v�gnar , f�r att han har efterstr�vat kompromisser i utskottet och funnit dem .
vad den fick fram var , med neil armstrongs , den ber�mde amerikanske astronautens , ord " ett j�ttespr�ng f�r m�nskligheten " , i det att de gick fr�n 350 gram till 50 gram i ett slag .
jag �r ledsen , ferber , jag bryr mig om f�rlorade arbetstillf�llen och den effekt som en s�dan f�rlust f�r .
en del av min grupp delar inte min �sikt p� ett antal punkter . det kommer ni strax att f� h�ra .
vad som skulle st�mma b�ttre �verens med medborgarnas f�rv�ntningar �r en �terst�lld j�mvikt i fr�ga om offentligt tillhandah�llande av tj�nster , genom att varje ny utvidgning till den kommersiella sf�ren f�rbinds med villkoret om en respekt f�r det grundl�ggande m�let om en h�llbar utveckling av det europeiska samh�llet .
privata operat�rer kommer att kunna dela ut brev till fyra g�nger den allm�nna avgiften .
i det t�nker man sig en minimal ytterligare �ppning av marknaden och en total os�kerhet om framtida �tg�rder kvarst�r , fast�n exemplet sverige borde lugna alla som tror att privatisering inneb�r att de samh�llsomfattande tj�nsterna f�rsvinner .
�ven om det steg som parlamentet nu vill ta �r alltf�r litet , s� b�r vi i vilket fall som helst se till att vi kan plocka upp tr�den igen om ett antal �r .
georg och markus , jag s�ger bara : n�r brevb�raren ringer p� d�rren en g�ng , eller kanske tv� , �r det inte europas sista sociala instans .
som v�rt utskotts f�redragande f�r tj�nster av allm�nt intresse r�der det f�r mig inget som helst tvivel om att vi kommer att bli tvungna att kritiskt granska den h�r utvecklingen .
mina spanska kolleger s�ger - och jag skulle g�rna vilja att kommission�ren talar om ifall de har r�tt - att spanien i full utstr�ckning har utf�rt direktivet fr�n 1997 , att andra inte har gjort n�gonting och att alla de d�r andra som inte har gjort n�gonting , nu vill ta ett j�ttesteg .
i v�rt fall har t.ex. ett land med en andel vilken ligger mycket under genomsnittsv�rdet naturligtvis inte n�got problem medan ett land med en betydande avvikelse upp�t kommer i en hoppl�s situation om �ven den gr�ns�verskridande posten avregleras enligt herr bolkesteins f�rslag .
vi i den h�r f�rsamlingen m�ste ge postmarknaden en chans .
fru talman ! det statliga monopolet p� posttj�nster inf�rdes inte utan anledning p� artonhundratalet .
kommissionens f�rslag om att avreglera posttj�nsterna har diskuterats intensivt �ver hela min valkrets , fr�n malin head till connemara och fr�n dublins utkanter till �arna .
just utifr�n de spanska erfarenheterna , vilka har n�mnts vid n�got tillf�lle , anser jag att parlamentets �ndringsf�rslag f�rb�ttrar kommissionens f�rslag eftersom det f�r in en m�ttlighet - strikt m�ttlighet - i �ppnings- och avregleringstakten .
fru talman ! arlette laguiller och jag sj�lv mots�tter oss alla former av inf�rande av privat kapital i postsektorn .
fru talman , kommission�r bolkestein , kolleger ! det verkar som om �mnet f�r dagen �r en l�ngdragen process : tv� steg fram�t , ett steg bak�t , s� l�ngsamt g�r vi fram�t i en av de viktigaste politiska fr�gorna med avseende p� fullbordandet av den inre marknaden , avreglering av postsektorn .
det �r anledningen till att jag p� nytt har lagt fram n�gra av de �ndringsf�rslag som vi diskuterade i utskottet och som vi kommer att r�sta om - s�rskilt ang�ende avregleringen av direktreklam .
det kommer att bli ett trefaldigt slag f�r storbritannien och ett trefaldigt slag s�rskilt f�r den brittiska landsbygden : ett slut p� den dagliga utdelningen och h�mtningen ; ett slut p� enhetliga priser - m�nniskor p� landsbygden kommer att betala mer f�r sin post ; och f�r det tredje och sista , ett slut p� v�rt omfattande och utm�rkta n�tverk av mindre postkontor p� landsbygden .
det �r verkligen en balanserad kompromiss , och jag hoppas att det kommer att antas av r�det .
det �r p� samma s�tt i den h�r debatten : det h�gst�mda talet om att bygga upp europa d�ljer illa �ngsligheten och konservatismen .
se var vi st�r i dag , mer �n tio �r senare .
om vi g�r f�r lite , f�r sent , kommer postsektorn som helhet att �ventyras .
v�rt f�rslag �r en noggrann balansg�ng , eftersom tillhandah�llare av samh�llsomfattande tj�nster kommer att beh�va tid f�r att �ndra strukturerna ytterligare , i syfte att bli flexiblare f�retag , s� att de kan anpassa sig till de nya marknadsf�rh�llandena .
i den andan kan jag godta de av era �ndringsf�rslag som inte �r orimliga och andra som med r�tta betonar fr�gor som samh�llsomfattande tj�nster som de till�mpas i medlemsstaterna , pr�vning av klagom�l samt n�tverket p� landsbygden .
f�r det andra kommer hela denna fr�ga att diskuteras i r�det ( industri / telekommunikation ) p� fredag .
vi f�rs�kte n� fram till en f�rlikning med kommissionen , vilket inte riktigt lyckades .
vi uppr�ttade kontakter med kommissionen , och vid det sista sammantr�det bekr�ftade kommissionen att den st�r fast vid sin st�ndpunkt , dvs. ett tullkvotsystem f�rvaltat enligt regeln " f�rst till kvarn " och en �verg�ng till tariff only �r 2006 .
detta f�rslag har redan godtagits av ecuador som �r v�rldens st�rsta bananproducent och en av dem som har lagt in en anm�lan till v�rldshandelsorganisationen .
jag tycker inte att det �ndringsf�rslag som vatanen ingivit i sista minuten underl�ttar saker och ting , varf�r jag uppmanar er , om ni lyssnar , till att fundera p� att dra tillbaka det .
jag vill d�rf�r h�r p�minna om att bananproduktionen inte �r en fr�mmande produktion i gemenskapen .
wto �r en upps�ttning regler .
d� kommer vi troligtvis att ha en annan maktposition och det visar sig d� �ven i bananbet�nkandet och i den m�ls�ttning som vi d� fastst�ller .
dessa olika l�nder har kunnat utveckla sin produktion p� grund av att vi erbjuder dem en marknad som vi i dag inte f� dra undan f�r dem .
avslutningsvis vill jag gratulera f�redraganden , dary , till det utm�rkta arbete han har utf�rt .
jag vill ocks� tacka ordf�randen f�r utskottet f�r jordbruk och landsbygdens utveckling , graefe zu baringdorf , f�r arbetet med att n� en kompromissl�sning med kommissionen .
det �r mycket or�ttvist .
v�lkomsth�lsning
herr talman ! jag tackar f�r st�det fr�n alla grupper .
( talmannen f�rklarade den gemensamma st�ndpunkten godk�nd ( efter dessa �ndringar ) . ) ( sammantr�det avbr�ts kl .
d�remot �r kommissionen beredd att godta �ndringsf�rslag 1 , 2 , 3 , 5 , 11 , 12 , 13 , 14 och 15 .
det godk�nner ocks� �ndringsf�rslagets f�rfattare .
bet�nkande ( a5-0376 / 2000 ) av theato f�r budgetkontrollutskottet om kommissionens meddelande om skydd av gemenskapernas ekonomiska intressen - bedr�geribek�mpning - f�r en gemensam �vergripande strategi ( kom ( 2000 ) 358 - c5-0578 / 2000 - 2000 / 2279 ( cos ) )
. ( el ) tyv�rr har r�det f�rkastat de flesta av europaparlamentets �ndringsf�rslag till skillnad fr�n kommissionen som har godtagit flera av dem .
med juridiska argument som t�ckmantel har vissa ledam�ter i europaparlamentet i realiteten f�rsvarat tobaksindustrin .
vi har ingen r�tt att diktera f�r andra vad de skall g�ra i sina l�nder utanf�r eu , och det �r inte heller s�rskilt klokt att exportera arbetstillf�llen fr�n eu till tredje land , d�r man helt enkelt kommer att framst�lla och s�lja produkterna och ta �ver v�ra nuvarande marknader .
s� mycket som en halv miljon m�nniskor i europa d�das av tobaken , och 85 procent av all lungcancer orsakas av r�kning .
herr talman ! jag r�stade f�r trakatellis bet�nkande i vilket det som vi vet avs�tts 79,1 miljoner euro f�r 2001-2002 , av vilka 8,5 till h�lsoupplysning , 31,1 till kampen mot cancer , 22,2 till f�rebyggande av aids , 11,4 till kampen mot narkotikaberoende , 4,4 till h�lso�vervakning och 1,3 till kampen mot sjukdomar till f�ljd av milj�f�rst�ring .
herr talman ! jag r�stade f�r detta direktiv om f�retag som f�r �vertagandebud .
det kan , d�rf�r , inte vara parlamentets m�l att undergr�va den europeiska konstmarknaden , och jag hoppas nu att medlemsstaterna och kommissionen kommer att kunna f�rsvara den gemensamma st�ndpunkten .
av dessa sk�l r�star de gruppl�sa nej till bet�nkandet .
dessutom kommer b�de unga och v�lrenommerade konstn�rer att lida av att den internationella handeln till f�ljd av en europeisk �verreglering kommer att utspela sig utanf�r europas gr�nser .
i allm�nhet �r t.ex. de finansiella medel som ansl�s till stabiliseringen av detta omr�de notoriskt otillr�ckliga .
situationen �r alarmerande .
bedragarna kommer att v�lja ut de l�nder som har det s�msta skyddet .
i corpus juris f�rutses det eventuella inr�ttandet av en oberoende europeisk �klagarmyndighet , med jurisdiktion f�r brott mot eu : s ekonomiska intressen som utf�rs b�de av ledam�ter och tj�nstem�n inom eu : s institutioner och av tredje part .
om jag i den processen kan skydda v�ra avs-l�nders intressen , s� �r det bra , men jag anser att det �r viktigt att vi skyddar och s�rjer f�r de europeiska medborgarnas v�lf�rd .
i darys bet�nkande �r man med fog orolig f�r s�v�l gemenskapens bananproducenter som avs-l�nderna .
jag kan �ven godta �ndringsf�rslag 28 , om en motsvarande best�mmelse l�ggs till om m�jligheten till en minskning .
enligt kommissionens uppfattning �r de tio �r som kr�vs i �ndringsf�rslag 11 och 13 f�r l�ng tid .
toppm�tet eu / usa
vi skulle vilja inrikta dessa toppm�ten , som �ger rum tv� g�nger om �ret , p� strategiska fr�gor som kan str�cka sig �ver flera toppm�ten .
avslutningsvis �r jag s�ker p� att vi kommer att ber�ra besluten nyligen i nice om den europeiska insatsstyrkan .
det viktigaste kommer att vara att vi g�r en konsolidering , att vi tar oss en noggrann titt p� hur de olika program ser ut som vi har initierats inom ramen f�r den transatlantiska dagordningen .
jag vet att kommissionen nu talar om att f�rnya delar av sin st�ndpunkt inf�r en ny runda , f�r att g�ra den flexiblare , och jag ser fram emot att f� veta vad det egentligen inneb�r i praktiken .
vi kan om�jligen acceptera att den enda l�sningen p� brott och v�ld skulle vara brott och v�ld .
det skulle vara ett n�je f�r oss att i den analysen innefatta en �versikt av det s�tt som de olika dialogerna har utvecklats p� .
vi b�r alltid f�rsvara den st�ndpunkten , utan att t�nka att vi genom att g�ra det p� n�got s�tt undergr�ver v�rt f�rh�llande till v�ra st�rsta v�nner och allierade .
min milit�ra karri�r var varken l�ng eller lysande , men jag l�rde mig att syftet med artilleriet var att bombardera infanteriet , det fientliga infanteriet om det var m�jligt .
f�r det andra , tj�nster avseende digitala produkter �r tj�nster och inte varuleverans .
i denna situation har kommissionen genomf�rt en studie om vad man kan g�ra , den vi behandlar h�r .
avslutningsvis vill vi s�ga att vi inte tycker om att se att kommissionen i b�rjan av sitt mandat fullkomligt l�mnar harmoniseringen av merv�rdesskatten d�rh�n och att parlamentet , �ven om det inser att det �r n�dv�ndigt att f�rl�nga giltighetstiden f�r g�llande lagstiftning , skall v�nta p� att kommissionen i mitten av sin mandatperiod och med euron redan i omlopp , skall l�gga fram ett nytt komplett och grundligt f�rslag i fr�gan .
i den bem�rkelsen v�lkomnar jag kommissionens tappra f�rs�k att finna ett s�tt att sluta det konkurrensgap som helt klart finns mellan e-aff�rer inom och utanf�r eu .
allteftersom t�gtrafiken byggs ut och erbjuder ett likv�rdigt alternativ , b�r man fr�mja det alternativet .
jag tror att det b�sta ur r�ttvisesynpunkt f�r de olika transportsektorerna , samt ur konkurrenssynpunkt , �r att vi g�r f�re och inf�r flygbr�nsleskatt i eu .
d�remot vet vi alla numera att en oreglerad konkurrens p� skatteomr�det �r en nackdel f�r alla .
d�remot m�ste en uppdelning ske av skatteint�kterna mellan medlemsstaterna p� grund av den stora sp�nnvidden p� satserna f�r merv�rdesskatt , precis som v�r f�redragande s� riktigt f�resl�r .
det kr�vs ett globalt syns�tt .
det skulle ocks� skapa st�rre r�ttvisa mellan olika transportslag .
jag kan , till exempel , inte f�rst� varf�r eurons inf�rande skulle kr�va en ytterligare eller ens n�gon samordning av merv�rdesskattesatser .
vi �r medvetna om v�ra riktv�rden : vid en skattesats p� mer �n 45 procent uppst�r i ett stort antal av v�ra medlemsstater ett budgetunderskott . riktv�rdena f�r usa �r andra .
jag skulle vilja uppmana kommissionen att ompr�va f�rslaget och att fundera p� en alternativ v�g .
samordna , harmonisera , betyder inte att likrikta .
herr talman ! det �r verkligen r�rande att lyssna till de �nglalika f�rsvarstalen f�r den elektroniska handeln , men det problem vi har h�r �r en reell konkurrensnackdel f�r v�ra europeiska f�retag , och vi m�ste r�tta till denna situation genom att fastst�lla vissa best�mda spelregler , s� att alla tj�nster som tillhandah�lls privatpersoner p� elektronisk v�g i europeiska unionen �r momsbelagda .
det �r just det vi vill skall ske med flygplanen !
vidare ligger det h�r f�rslaget , i mina �gon , i linje med de principer som man har kommit �verens om i ekofin-r�det , vilka i sin tur ligger i linje med de principer som man enades om vid oecd : s konferens i ottawa .
n�r flygbiljetterna �r 42 procent billigare i dag �n f�r tio �r sedan , �r det uppenbart att felaktiga prissignaler s�nds ut .
allm�nheten f�rtj�nar n�gonting b�ttre .
jag delar inte den uppfattningen .
herr talman ! jag anser att tanken p� en ensidig upps�ttning best�mmelser f�r beskattning av br�nsle f�r luftfartyg i eu inte alls �r �ndam�lsenlig , mot bakgrund av att vi globalt fortfarande �r underst�llda chicagokonventionen fr�n 1944 , som undantar flygfotogen fr�n beskattning internationellt .
den skapar r�ttss�kerhet f�r varje enskild sparare och medborgare .
sedan kommissionen presenterade f�rslaget den 7 juni i �r har den saken f�tt mycket uppm�rksamhet de senaste m�naderna .
det �r en f�rdel att det finns ett klart och objektivt kriterium , n�mligen den medlemsstat d�r konsumenten bor .
det �r en f�renklings�tg�rd som reglerar utbytet av information om momsregistreringsnummer i den elektroniska handeln mellan medlemsstaterna , och vi kommer att l�gga f�rslaget p� minnet i v�rt fortsatta arbete i parlamentet och r�det .
dessa diskussioner kommer emellertid att bli mycket sv�ra med tanke p� att man under den f�reg�ende f�rsamlingen inte n�dde fram till n�got beslut om m�jligheten att inf�ra beskattning av br�nsle f�r luftfartyg .
denna olycka , som var en i raden av m�nga andra , v�ckte de ber�rda befolkningarnas , liksom den �vriga allm�nhetens , vrede och missmod inf�r sj�fartens ogenomtr�nglighet och sv�righeter att anpassa sig till g�llande best�mmelser f�r att undvika denna typ av problem .
det andra m�let �r att vid olyckor f�renkla och skynda p� en detaljerad informationsf�rmedling om farlig eller f�rorenande last och tvinga fartygen och myndigheterna att meddela uppgifterna p� elektronisk v�g .
betr�ffande ansvarighetsfr�gan : den m�ste vi granska ing�ende .
n�r det g�ller f�rdskrivaren skall vi s�ga att internationella sj�fartsorganisationen planerar ett obligatorium av denna typ f�r de fartyg som seglar p� nationella rutter fr�n och med juli 2008 , men vi vill tidigarel�gga detta datum .
herr talman ! jag skulle i min tur vilka tacka palacio f�r hennes uttalande .
fr�ga nr 33 fr�n ( h-0873 / 00 ) :
�r det allts� godtagbart att fordon kan stoppas vi gr�nsen till en angr�nsande medlemsstat , trots att de uppfyller alla krav i det egna landets lagstiftning ?
de bidrar s�ledes inte alls till infrastrukturkostnaderna f�r v�gar i storbritannien och betalar samtidigt l�gre fordonsskatter i hemlandet .
. ( en ) jag har ingen m�jlighet att ge er exakta siffror om m�ngden importerat k�tt fr�n tredje land , men jag kan s�ga att den importen styrs av de l�mpliga f�reskrifterna och att �verv�ganden om livsmedelss�kerhet ligger till grund f�r den lagstiftningen .
herr talman ! judarna �r profeternas och de troendes fiender .
s� jag upprepar : vi kommer att diskutera fr�gan med de palestinska myndigheterna .
koncentrationsf�rordningen erbjuder ingen r�ttslig grund f�r att beakta p�st�enden om brott mot de m�nskliga r�ttigheterna , och kommissionen har d�rf�r inga befogenheter att unders�ka s�dana p�st�dda brott i detta sammanhang .
omv�nt st�r andra medel till medlemsstaternas och europeiska unionens f�rfogande f�r att hantera fr�gor som r�r de m�nskliga r�ttigheterna .
dessutom kommer kommissionen , om den inte , inom ramen f�r f�rfarandet enligt handelshinderf�rordningen , n�r en f�rhandlingsl�sning med korea som �r tillfredsst�llande f�r europeiska unionen , att rapportera till r�det senast den f�rsta maj 2001 och f�resl� att fallet tas till wto , i syfte att s�ka motmedel mot illojala koreanska metoder .
vi f�r inte heller gl�mma att valdivielso de cu� fr�gade er om kommissionen trodde att denna varvsindustri hade �verlevt i europeiska unionen utan de st�d den har f�tt .
syssels�ttningsfr�gan har f�tt en s�rskild uppm�rksamhet .
ang�ende : f�rslaget om att avskaffa importtullarna f�r samtliga varor utom vapen n�jer sig kommissionen med att detta dramatiska f�rslag - som mycket v�l kan f� �desdigra konsekvenser f�r de redan h�rt ansatta sockerbetsodlarna i europeiska unionen - skulle antas utan att det direktvalda europaparlamentet ombeds yttra sig ?
n�r det g�ller fr�gan som st�lldes av glenys kinnock , huruvida detta initiativ �r f�renligt med avtalet fr�n cotonou , skulle jag �n en g�ng vilja s�ga att kommissionen till fullo har respekterat s�v�l andan som ordalydelsen i avtalets best�mmelser om information till och samr�d med avs-l�nderna .
det st�mmer att sockerpriset i europeiska unionen i dag �r tre g�nger h�gre �n p� v�rldsmarknaden , vilket verkligen st�ller till med problem .
betr�ffande fr�gan huruvida det �r en taktisk gest som �r avsedd att locka till sig fav�rer fr�n de minst utvecklade l�nderna inom ramen f�r en f�rhandlingsrunda , vill jag genast klarg�ra att s� inte �r fallet .
en av de fyra organisationerna �r ecpat , vars st�dber�ttigade �tg�rder inom detta omr�de under 2001 helt omfattas av denna ans�kan .
herr talman , �rade kommission�r liikanen ! vi kommer sent i kv�ll att diskutera direktivet om digitalt inneh�ll .
en ny artikel i f�rdraget m�jligg�r en eventuell utvidgning av eg-domstolens befogenheter i det h�r avseendet .
jag skulle vilja f�rs�kras om att kommissionen kommer att �verv�ga f�rdelarna med ett s�dant tillv�gag�ngss�tt mycket noga , eftersom jag misst�nker att en f�r�kning av jurisdiktionsomr�den i slut�ndan kan splittra v�ra r�ttssystem .
vilka �tg�rder t�nker kommissionen vidta f�r att se till att de medlemsstater som �nnu inte gjort det utser domstolar f�r gemenskapsvarum�rken ?
jag tackar herr berenguer fuster f�r att han framst�ller en s� stark beg�ran till kommissionen .
herr kommission�r ! jag m�ste erk�nna att ni inte har informerat mig eller snarare att ni inte har sagt n�got nytt som jag inte redan visste eftersom ni sedan ett �r tillbaka har detta klagom�l hos kommissionen .
tack f�r svaret , herr kommission�r .
det r�r sig i det fallet om en brittisk examen .
fr�ga nr 49 fr�n ( h-0912 / 00 ) :
man letar som b�st efter andra l�nsammare fartyg och transportf�retag i st�llet f�r dem som nu slutar , med avsikten att f�rena person- och frakttrafiken .
herr talman ! jag v�lkomnar detta initiativ fr�n kommissionen .
det �r d�rf�r n�dv�ndigt att f�rkorta programmets till�mpningsperiod , vilket g�r att programmet kan f� mycket st�rre effekt , tack vare att mer pengar skjuts till under en kortare tidsrymd .
jag skulle vilja veta vad som kommer att ligga i ordet " inneh�ll " .
f�rmedlingen av digital information saknar gr�nser av tidigare slag .
europeiska folkpartiets grupp och europademokrater kommer h�r att ta fasta p� f�rslagen - och det tackar jag gill f�r - , �ven vi kommer att r�sta f�r ett h�jt bidrag och jag hoppas att denna �verenskommelse med europeiska liberala , demokratiska och reformistiska partiets grupp och andra grupper skall h�lla , att vi verkligen kommer att k�mpa f�r det , att dessa budgetposter verkligen kommer att ut�kas , s� som vi har f�reslagit .
faktum �r att den lovordade kulturella och spr�kliga m�ngfalden i europa ofta �r ett hinder , framf�r allt f�r den gemensamma marknaden .
det �r s�ledes ett mycket viktigt program och ett mycket viktigt bet�nkande , och f�r detta vill jag gratulera kommissionen , kommission�r liikanen och fru gill .
vi m�ste se till att det finns en milj� som kan underl�tta dessa f�r�ndringar i europa .
de �terst�ende 11 �r inte direkt f�renliga med m�len i det h�r specifika programmet , eller s� skulle de str�cka programmets mandat bortanf�r gr�nsen f�r vad som kan uppn�s med de ekonomiska medel som �r f�rknippade med det .
jag skulle emellertid vilja uppmana ppe-de-gruppen till att i vilket fall som helst inte st� i v�gen f�r att diskussionen om saken �ger rum nu i kv�ll .
( �terf�rvisning av bet�nkandet till utskottet f�rkastades . )
subsidiaritetsprincipen - det kommer snart att visa sig i debatten - �r ett viktigt element . �ven den vill utskottet f�r milj� ta h�nsyn till .
nu n�r omgivningsbullret har stigit kraftigt , inte minst till f�ljd av den �kade r�rligheten , s� har ocks� antalet m�nniskor som konfronteras med det v�xt starkt .
f�redraganden har n�mnt en mycket h�gre procentsats , och faktum �r att omgivningsbuller �r ett stort och allvarligt milj�problem .
f�redraganden �r mycket kreativ i sina f�rslag om ramdirektiv och f�ljddirektiv samt f�rslaget om att g�ra bullerkartor tillg�ngliga f�r allm�nheten .
det st�r ett antal bra och viktiga saker i det h�r direktivet , harmoniseringen , bruket av gemensamma bullerm�tt och parametrar , programvara och liknande saker .
i spanien och i m�nga medelhavsl�nder �r den normala dagsl�ngden ganska mycket senare �n klockan 19.00 som detta direktiv anger .
vi m�ste f�lja den v�gen , men f�redraganden nuvarande f�rslag g�r f�r tillf�llet f�r l�ngt i den riktningen .
f�r det f�rsta m�ste vi ha ett ramdirektiv d�r m�tmetoderna och handlingsplanerna fastst�lls , och en standardisering av politiken p� det omr�det m�ste skapas .
jag skulle vilja veta vilken slutsatsen egentligen var .
vi kommer att �verv�ga vilka dessa standarder beh�ver vara s� snart vi har ett underlag fr�n strategiska bullerkartor .
kommissionen kan godta �ndringsf�rslagen 1 till 3 , 14 , 18 , 27 , 30 , 34 , 35 och 43 .
man kan f�rst� att alginatbehandlingen riskerar att vilseleda konsumenten eftersom den f� en produkt att se " f�rskare " ut �n den egentligen �r .
jag tror att det vore bra f�r folkh�lsan , samtidigt som det inte medf�r n�gra som helst skador f�r industrin .
f�r det andra , var finns industrins beredskap att stiga fram och godta att n�gra av de m�nga tillsatser som vi anv�nder kan tas bort ?
officiell kontroll p� djurfoderomr�det
under trepartsm�tet framgick det tydligt att r�det inte skulle ge efter p� den punkten .
hur kan man dock ge garantier n�r inga kontroller utf�rs ?
vi m�ste akta oss f�r att anv�nda ett tillv�gg�ngss�tt uppifr�n och ner f�r vad som bara kan vara ett initiativ nerifr�n och upp .
programmet f�r f�rnyelse av sm� st�der och byar �r en integrerad del av landsbygdens utveckling .
begreppet h�llbar utveckling , s�rskilt n�r det g�ller st�derna , �r inte enbart begr�nsad och kan inte enbart begr�nsas till milj�aspekten , utan har �ven sociala och ekonomiska aspekter .
b�ttre kunskap och ny teknik ger m�jligheter till b�ttre milj� i europas st�der .
det kommer att g�ra det m�jligt f�r och uppmuntra st�der runtom i europa och annorst�des att m�tas och l�ra av varandras erfarenheter , hj�lpa dem att angripa problem och utmaningar p� milj�omr�det och att arbeta i riktning mot en h�llbar utveckling .
den andra fr�gan g�ller kommitt�f�rfarandet .
. ( fr ) herr talman , herr kommission�r , k�ra kolleger ! det �r visserligen sent p� kv�llen som vi behandlar denna beryktade f�rsiktighetsprincip .
texten fr�n utskottet f�r milj� �r resultatet av ett st�ndigt s�kande efter en kompromiss , eller snarare en j�mvikt mellan maximalistiska och minimalistiska uppfattningar , som har uttryckts under v�ra debatter och som b�da utmynnar i �verdrifter .
vi m�ste s�kerst�lla att det h�r bet�nkandet �terspeglar allm�nhetens krav p� en h�g skyddsniv� f�r h�lsa och milj� .
f�rsiktighet �r n�dv�ndig i situationer d�r riskerna k�nda .
det gl�der mig f�ljaktligen att se att det slutliga bet�nkandet speglar behovet av att utveckla begreppet ytterligare .
d�r f�resl�s att omv�nd bevisb�rda skall till�mpas vad g�ller produkter utan f�rhandsgodk�nnande , det vill s�ga att producenten skall bevisa att produkten �r s�ker och inte �verl�ta riskerna och kostnaden p� konsumenterna .
som alla vet genomsyras livet av risker och tveksamheter .
� andra sidan anv�nds det �ven av europeiska unionen p� ett ganska otydligt och till och med irrationellt s�tt .
men det finns fler exempel �n galna ko-sjukan , exempel som kanske inte �r lika spektakul�ra , men d�r det �r lika viktigt att vi fattar beslut .
en analys av f�rdelarna och nackdelarna �r en absurd id� , n�r man t�nker p� vad som �r syftet med f�rsiktighetsprincipen , n�mligen att kunna reagera p� en produkt redan innan man k�nner till alla f�rdelar och nackdelar .
f�rsiktighetsprincipen diskuterades �ven vid toppm�tet i nice , som tog notis om en resolution som antagits av r�det ( allm�nna fr�gor ) .
det �r viktigt att betona att det �r upp till beslutsfattarna att best�mma skyddsniv�n .
i detta uttalande f�rd�mer vi kraftfullt eta : s brott i spanien , och europeiska unionens institutioner uppmanas att vidta effektivare �tg�rder f�r att bek�mpa terrorismen .
( livliga och ih�llande appl�der )
valda icke-nationalistiska politiker m�rdas liksom f�retagare , journalister , anst�llda i den allm�nna ordningsmakten eller bara enskilda som p� n�got s�tt har uttryckt sig emot det tv�ngsm�ssiga sj�lvst�ndighetsprojektet .
jag �r dock givetvis h�nvisad till sessionstj�nstens f�rarbete .
vi skall �terl�mna faderskapet till er .
f�re omr�stningen om �ndringsf�rslag 51
( parlamentet antog resolutionen . )
att stora schweiziska milj�organisationer har l�tit sig �vertalas med argumentet att inkomsterna fr�n avgifter skall g� till en utbyggnad av j�rnv�garna �vertygar mig inte alls .
vi gl�der oss �t att detta h�danefter �r erk�nt .
i luxemburg f�r p� sin h�jd tekniska tj�nster som tryckerier och �vers�ttningstj�nsten finnas kvar .
budgeten f�r 2001 bygger i stor utstr�ckning p� en kompromiss mellan parlamentet , r�det och kommissionen , som vi st�ller oss bakom .
d�rmed , och f�rvisso mycket sent , erk�nner europeiska unionen s�ledes h�danefter hur viktig en omfattande hj�lp till den sv�rt �rrade jugoslaviska republiken �r med respekt f�r dess gr�nser .
detta �r en p�fallande svag slutsats .
genom att den europeiska marknaden stegvis avregleras , kan posttj�nsterna effektiviseras och servicen till kunderna h�jas .
. ( fr ) hur kommer postsektorn att ta sig ur denna period d� mots�gelser och tvister har kommit f�r att ofta nog st�dja tekniska f�rsvarstal som utarbetats inom ramen f�r sektorns �ppnande f�r konkurrens ?
pris- och viktgr�nserna fastst�lls p� ett f�rnuftigt s�tt , det vill s�ga att upp till 150 gram f�rbeh�lls de samh�llsomfattande posttj�nsterna , liksom �ven en prisgr�ns som uppg�r till fyra g�nger den allm�nna tariffen .
- ( pt ) kommissionens f�rslag f�r postsektorn inneb�r en avregleringsvilja utan gr�nser , och �r en attack p� en viktig offentlig service och p� de f�retag och de anst�llda som utg�r dem .
europaparlamentet ger allts� kommissionen en stark signal om sina reservationer inf�r en totalt avreglerad postmarknad .
jag anser inte att europeiska unionens pengar skall anv�ndas p� detta s�tt !
vi har inte f�r avsikt att vare sig gynna de stora hajarna i bananbranschen eller de mellanstora hajarna i det omr�de som skyddas av europa .
h�rmed tillhandah�lls i europakonventionen om skydd av m�nskliga r�ttigheter och grundl�ggande friheter en ram f�r begr�nsning av inneh�ll i syfte att skydda anv�ndare .
. ( fr ) programmet econtent syftar till att uppmuntra utveckling och utnyttjande av europeiskt digitalt inneh�ll i de globala n�ten samt fr�mja spr�klig m�ngfald i informationssamh�llet .
n�r det g�ller det digitala , inneb�r det spr�kliga uttrycksmedlet samtidigt ett konkurrens�vertag , ett tankes�tt och en r�ttslig �terverkan som gynnar dem som har det som modersm�l .
� andra sidan hyser jag hopp inf�r den regeringskonferens som skall ske �r 2004 , som �r det enda som jag tycker �r positivt fr�n nice , s� att denna en g�ng f�r alla beaktar f�rdelning och distribution av kompetenser mellan europeiska unionen och l�ndernas regeringar .
. ( fr ) europeiska r�det i nice hade en positiv sida : genom att visa upp en ny r�stviktning och en ny f�rdelning av de europeiska parlamentsledam�terna som b�dadera omfattar kandidatl�nderna fr�n �steuropa har det just gett dessa ett tydligt tecken p� sin vilja att ta emot dem p� kort sikt .
trots en l�tt h�jning av tr�skeln f�r kvalificerad majoritet , vars omfattning m�ste kontrolleras , borde detta breddande inneb�ra att klyftan ytterligare kommer att �ka mellan de europeiska institutionerna och de nationella demokratierna .
flera medlemmar av europaparlamentet har uttalat sig mycket kraftfullt f�r en utvidgning av dagordningen .
vi har �nnu n�gra m�nader p� oss fram till slutet av 2003 f�r att r�dda det europeiska projektet .
trots de framg�ngsrika initiativ som togs p� detta omr�de under toppm�tet i nice , uttrycker resolutionen missn�je med den nya utvidgningen av de kvalificerade majoritetsbeslutens r�ckvidd .
tv�rtom : de europeiska medborgarna och deras parlament upplever nu ett steg tillbaka fr�n amsterdam .
faktum �r att inget toppm�te hittills har tvingats ta itu med en s� stor utvidgning som denna .
inga steg tas f�r att g�ra eu mer demokratiskt eller �ka de nationella parlamentens makt .
vi pension�rer reser ofta och om sanningen skall fram �r det anstr�ngande att resa med t�g eller bil : f�r oss �r flyget en dr�m som f�rverkligas .
" d� g�r jag till fots .
det �r ett f�rs�k som �r v�rt att st�dja , eftersom klyftan mellan de mest utvecklade och de minst gynnade regionerna �r mycket st�rre n�r det g�ller den tekniska utvecklingen �n f�r bruttonationalprodukten .
herr talman ! l�t mig i en mycket positiv anda kommentera markovs bet�nkande och gratulera honom till att ha lagt fram ett s� konstruktivt bet�nkande f�r kammaren .
d�rf�r b�r inte innovationsfaktorer nedv�rderas av n�gon , hur obetydliga de �n m� vara , som denna .
just den tekniken ger dem nu ett redskap f�r att ta igen denna eftersl�pning under f�ruts�ttning att de ekonomiska akt�rerna i regionerna �ven �r i st�nd att anv�nda de innovativa �tg�rderna f�r att utnyttja den m�jligheten .
i konsekvensens namn m�ste denna uppmaning naturligtvis �tf�ljas av en begr�nsning av den besv�rliga byr�kratin , herr kommission�r , p� alla niv�er , n�r det g�ller ig�ngs�ttande och genomf�rande av programmen .
det var s�rskilt positivt att i synnerhet kvinnorna fick engagera sig i fr�gan om den nya tekniken .
f�rutom detta tas , som en konsekvens av v�r komplexa institutionalisering , beslut p� gemenskapsniv� ofr�nkomligen l�ngsamt . d�rf�r �r det inte f�rv�nande att vi finner att vi inte ens kunnat g�ra av med den budget som f�rutsetts f�r innevarande �r f�r innovativa �tg�rder i den regionala politiken och det �r en politisk oansvarighet .
i samband med de prioriterade teman som valts och som jag personligen ville l�gga fram inf�r utskottet f�r regionalpolitik den 11 september , skulle jag vilja upprepa att dessa innovativa �tg�rder framf�r allt �r ett instrument f�r regional utveckling .
vi har dessutom tagit upp vissa aspekter f�r att g�ra det m�jligt f�r sm� och medelstora f�retag att finna l�sningar p� behoven n�r det g�ller datakunskaper och personalen .
jag m�ste liksom ni n�ja mig med de medel som planerats i riktlinjerna fr�n berlin och paketet i agenda 2000 .
enligt kommissionens rapport har sydkorea i �rets best�llningar hittills kammat hem mer �n 40 procent av alla best�llningar p� fartygsbyggen p� land , och det tack vare krediter fr�n sydkoreanska banker som till viss del �gs av staten , tack vare statliga garantier som motsvarar subventioner .
jag hoppas att den valda tidpunkten f�r presentationen av denna rapport f�r parlamentet inte var ett knep f�r att uppmuntra oss till att ta bort denna punkt fr�n f�redragningslistan .
vi har ocks� framf�r allt noterat r�dets slutsatser fr�n den 5 december . ett r�d som har accepterat att skydda framtiden genom att visa fasthet gentemot sydkorea och genom att inte st�nga d�rren f�r m�jligheten att �teruppr�tta st�det till varvsindustrin i maj n�r det g�ller best�mda marknadssegment som kraftigt drabbats av den koreanska konkurrensen .
jag anser att det �r s� att vi i europa lider av en illojal konkurrens eftersom man i korea f�rst och fr�mst betalar mycket l�ga l�ner , i kombination med hemska arbetsvillkor f�r de koreanska arbetstagarna , och under dessa villkor kan de europeiska arbetstagarna inte p� n�got s�tt konkurrera med dem .
med denna form av bidrag , vilken �r �ppen f�r insyn , �r det inte lockande f�r europeiska varv att till�mpa olika rabatterings- och marknadsf�ringsmetoder som inte �r f�renliga med marknaden .
d�r �r nu det som tidigare var skeppsvarv ett konserthus och sj�fartsmuseum , etc . tidigare arbetade 4000 personer p� varven men nu arbetar tv� vaktm�stare p� varje st�lle , och det �r vad som sker i de europeiska l�nderna .
herr talman ! jag skulle vilja inleda med att gratulera langen f�r kvaliteten i hans bet�nkande .
som ett resultat av detta misslyckande formulerade industrin ett klagom�l i oktober i �r , i enlighet med f�rordningen om handelshinder ( tbr ) , och kommission�r lamy meddelade den 4 december kommissionens beslut att inleda en unders�kning .
detta f�rslag kommer att l�ggas fram om det inte g�r att �stadkomma ett tillfredsst�llande avtal med korea under loppet av unders�kningsf�rfarandet enligt f�rordningen om handelshinder .
han var en arbetare och som de som var med oss i g�r n�r vi delade ut sacharovpriset var han en anonym medborgare som tj�nade det demokratiska system spanjorerna har valt .
det var en g�ng en engelsk atomub�t som hette tireless .
ledam�ter , det handlar inte om att oroa .
i b�da beg�r vi att kommissionen skall utr�na m�jligheterna i de nuvarande f�rdragen f�r att ta reda p� vilka m�jligheter den har att bidra i denna fr�ga .
s�ledes har vi de h�r m�naderna deltagit i en rad av galenskaper .
hon beklagar att hon inte kan vara h�r och besvara fr�gorna personligen , men hon sitter i sammantr�de i bryssel och f�rbereder n�sta veckas viktiga ministerm�te om klimatf�r�ndringar .
som svar p� om det finns en interventionsplan f�r gibraltaromr�det och gibraltars hamn , har de brittiska myndigheterna informerat kommissionen om sin s�kerhetsplan f�r allm�nheten i gibraltar , k�nd under namnet " gibpubsafe " , som allts� �r interventionsplanen f�r gibraltar .
den f�rsta punkten jag vill ta upp �r att reparationerna av denna ub�ts kylsystem redan p�g�r .
problemet med ub�ten m�ste l�sas i lugn och ro och genom ett fullst�ndigt samarbete mellan alla ber�rda , beh�riga myndigheter .
kanske �r h�ndelsen allvarlig och kanske �r den det inte .
han beklagar sig �ver det . vi gl�der oss �t det :
denna situation kan inte p� n�got s�tt vara en bilateral fr�ga mellan tv� stater som tillh�r en politisk union .
gibraltars och s�dra spaniens befolkningars intressen �r identiska i detta avseende .
den spanska regeringen har hela tiden haft en inst�llning som grundar sig i tv� utg�ngspunkter : behovet av en �ppen information , med grund i tekniska och vetenskapliga kriterier f�r att bed�ma vidden av reparationen och dess riskpotential och ocks� det att varje slags beslut , vare sig om en reparation i gibraltar eller om en f�rflyttning till en bas i storbritannien skulle tas i enlighet med rigor�sa tekniska kriterier .
b5-0901 / 2000 fr�n sylla m.fl. , f�r gue / ngl-gruppen ;
det riktiga sk�let �r inte heller jubileet , utan snarare den n�dsituation som fn : s flyktingkommissariat befinner sig i .
detta �r emellertid inte tillr�ckligt , vi b�r m�lmedvetet st�dja unhcr politiskt och ekonomiskt f�r att garantera b�ttre prognoser , flexibilitet och geografisk balans .
alla som bes�kte den senaste utst�llningen i europaparlamentet och som studerade bilderna och texten som handlade om unhcr : s arbete i v�rlden just nu , tror jag skulle h�lla med om att det var en av de sorgligaste utst�llningar vi n�gonsin haft oturen att se i v�rt parlament .
dessa m�ten b�r hj�lpa kommissionen att tillhandah�lla en mer f�ruts�gbar och �ppen finansiering , som unhcr beg�r och har efterlyst sedan l�nge , samtidigt som den kan hj�lpa unhcr att bist� de beh�vande p� ett b�ttre s�tt .
b5-0902 / 2000 fr�n morgantini och frahm , f�r gue / ngl-gruppen ;
det �r ett andra problem .
den nya politiska ledningen i serbien m�ste agera p� ett s�dant s�tt , och detta vill jag po�ngtera , herr talman , s� att den f�rre presidenten och diktatorn milosevic , tillsammans med sina medf�rbrytare , kan f�ras till den internationella krigsf�rbrytartribunalen i haag .
vi f�rv�ntar oss antingen en klar amnestilag p� kort sikt med konkreta detaljer , eller , och helst i kombination , ett konkret datum f�r frigivning av de politiska f�ngarna .
det �r s� mycket som f�r�ndrats sedan i h�stas : de nya myndigheterna i belgrad har agerat snabbt , t.ex. f�r att �terst�lla sina internationella kontakter ; de har agerat snabbt f�r att g�ra det m�jligt f�r f�rbundsrepubliken jugoslavien att inta sin plats i f�renta nationerna och �ven i osse .
b5-0911 / 2000 fr�n grosset�te , f�r ppe-de-gruppen ;
m�nskliga r�ttigheter i tunisien- b5-0905 / 2000 fr�n boudjenah m.fl. , f�r gue / ngl-gruppen ;
och vid ett tillf�lle fick general pinochet f�r sig att komma till europa , och fr�n det att han satte f�tterna p� europeisk mark best�mde sig de europeiska r�ttsliga myndigheterna f�r att f�rs�ka uppn� att general pinochet skulle st� till svars f�r sina handlingar .
jag bekr�ftar ocks� st�det fr�n min grupp f�r �ndringsf�rslaget fr�n gruppen europeiska f�renade v�nstern / nordisk gr�n v�nster om milit�r inblandning i processen .
ett fredligt och demokratiskt genomf�rande av politiska m�l �r inte bara ett medel f�r att uppn� ett m�l - det �r inneboende i alla v�rdefulla m�l .
s� l�nge situationen �r s�dan , kan landet inte komma i fr�ga f�r medlemskapsf�rhandlingar med europeiska unionen .
jag �r glad �ver det eftersom jag anser att n�r det inte �r en smakl�s l�tsad situation , �r hungerstrejken ett sj�lvmordsbeteende som mina personliga �vertygelser hindrar mig fr�n att uppmuntra .
vissa , s�som b�chir habib , �r i ett kritiskt tillst�nd .
trots att n�gra pass har �terl�mnats , �ven om president ben ali p� �rsdagen av sitt makttilltr�de h�ll ett tal om pressfrihet och f�rb�ttrade f�ngelsevillkor , konstaterar vi en allvarlig f�rs�mring av situationen f�r m�nskliga r�ttigheter i tunisien .
fortfarande �r minst 1 000 personer f�ngslade f�r sina �sikters skull .
den unge studenten b�chir habid hungerstrejkar sedan den 18 oktober .
jag deltog i �verl�mnandet av makten i f�rbundet f�r m�nskliga r�ttigheter en vecka innan det f�rsattes i konkurs .
( talmannen avbr�t talaren . )
man gjorde offentliga uttalanden efter dessa evenemang , d� man beklagade anv�ndningen av v�ld och st�dde �tg�rder f�r att st�lla de ansvariga inf�r r�tta .
p� det finansiella omr�det , och detta har direkt att g�ra med det som ledamoten tog upp - och det �r ett omr�de d�r vi har f�tt en viss erfarenhet fr�n andra l�nder , �r kommissionens f�retr�dare i f�rd med att trappa upp sina anstr�ngningar f�r att inom kort kunna starta tv� program : ett till st�d f�r journalister och det andra till st�d f�r icke-statliga organisationer .
att forts�tta denna politik kan bara leda till ett blodbad , liknande det som har intr�ffat i andra l�nder .
vi f�r �nska att de har mod att anta utmaningen , och vi f�r inte spara p� n�gon anstr�ngning f�r att hj�lpa dem .
f�r att dessa verkligen skall leda till att l�sa upp den nuvarande situationen �r det n�dv�ndigt att f�rst skapa villkor f�r att s�dana val skall kunna h�llas under civil fred och f�rsoning .
ouatara har inte ivoriansk nationalitet och det �r absolut normalt , s�som det skulle vara i var och en av v�ra stater att elfenbenskusten avl�gsnar fr�n nationellt ansvar dem som inte har ivorianskt medborgarskap .
under debatten om den brittiska ub�ten i gibraltar sade ni att den allm�nna s�kerhetsplanen f�r gibraltar skulle finnas tillg�nglig f�r kollegerna i kammaren .
herr talman ! jag f�ljer kollegan wurtz exempel och drar formellt tillbaka v�rt resolutionsf�rslag .
jag inser att detta kommer att ge upphov till debatt .
jag uppfattar ert inl�gg som en uppmaning till �kad arbetsiver .
vi vet mycket v�l att h�lsan inte �r en g�va som varar i evighet .
i bakgrunden st�r fn : s internationella �r f�r �ldre och det har varit av st�rsta vikt att man p� olika h�ll f�ster uppm�rksamhet vid hur de �ldres situation utvecklas i framtiden , till exempel i de l�nder som h�r till europeiska unionen .
p� den tiden var detta undantag , d� de flesta m�nniskor avled p� grund av sv�ra f�rh�llanden vid en relativt l�g �lder .
europeiska institutioner har knappt n�gra befogenheter p� detta politiska omr�de .
m�nniskor beh�ver varandras omsorg och uppm�rksamhet , de �r involverade i varandra .
�ren g�r . de anst�llda blir sjuka p� grund av arbetet , de betalar sina pensionsavgifter , sina sjukf�rs�kringsavgifter .
de m�nga fallen av f�rtidspensionering och de varierande gr�nserna f�r pensionering f�ruts�tter dock ett enormt arbete f�r omv�rdering av dessa politikomr�den vilka inte alla rymmer social medk�nsla .
detta p�minner mig om diskussionen p� 1960-talet , d� det handlade om att h�lla oss kvinnor borta fr�n arbetsplatserna .
jag gratulerar v�r f�redragande . �ven jag vill inleda med ett konstaterande som var och en utan sv�righet kan inst�mma i : europa �r med tanke p� �lderspyramiden en �ldrande kontinent .
som medlem av den visserligen inte officiella men faktiskt existerande fredagsklubben tillh�r jag liksom ni den skara av ledam�ter som �r n�rvarande �ven denna dag , och jag hoppas att vi kommer att lyckas med det �ven n�sta �r .
den som n�jer sig med att vara en genomsnittsm�nniska kommer aldrig att ge sig in p� det �ventyr som det inneb�r att leva som en engagerad m�nniska .
det �r viktigt att bedriva en konkret politik och genomf�ra s�rskilda program f�r olika kategorier av �ldre personer .
vi st�r helt visst inf�r v�ldiga utmaningar .
alla kan eller skall inte frivilligt sluta att yrkesarbeta .
( skratt och appl�der )
det vore d�rf�r l�mpligt att fastst�lla tidpunkten f�r f�rordningens ikrafttr�dande till den dag d� genomf�randef�rordningen antagits , f�r att de anslag som �r tillg�ngliga f�r �r 2001 inte skall g� f�rlorade .
f�r det f�rsta b�r vi titta p� jordbruksprodukterna ur h�lsosynpunkt : mer frukt , mer mj�lk och s� vidare .
vi vill f�rbli friska och n�ringsmedel �r helt enkelt grunden till ett sunt liv .
av denna anledning �r det n�dv�ndigt med �tg�rder f�r information och marknadsf�ring finansierade av europeiska unionen och medlemsstaterna , b�de f�r att bidra till att �teruppr�tta det skamfilade rykte jordbruket f�tt hos konsumenterna och f�r att i �vrigt f� erk�nnande f�r den utm�rkta kvaliteten hos den �verv�gande delen av v�ra jordbruksprodukter .
eller om man talar om att vi har ett underskott n�r det g�ller proteinf�rs�rjning .
det kan inte rimligen vara skattebetalarnas och unionens sak att finansiera reklamkampanjer till exempel f�r att man skall k�pa tulpaner eller �ta mera �pplen .
utgifterna under det senaste programmet sj�nk faktiskt mellan 1997 och 1998 .
mulder har r�tt n�r han s�ger att den europeiska jordbrukspolitiken �r konstruerad inte bara f�r mat men i det sociala syftet att beh�lla h�gsta m�jliga antal m�nniskor p� landsbygden .
den sista gruppen �ndringsf�rslag som kommissionen inte kan acceptera g�ller �ndringar , som inte st�r i samklang med sj�lva f�rslaget , som skulle kunna f� o�nskade f�ljder och i vilka f�rvaltningsrutiner f�resl�s , som inte har sin motsvarighet i sedvanlig praxis .
f�r det �r faktiskt riktigt att det �r n�dv�ndigt , men ocks� ber�ttigat , att g�ra reklam f�r den europeiska jordbruksmodellen .
redan den helige benedikt uppmanade sina munkar att konsumera en halv tunna vin till varje m�ltid f�r att g�ra dem mera kvickt�nkta och f�r att f�rb�ttra deras matsm�ltning .
jag tycker verkligen att detta �r alldeles f�rskr�ckligt , det strider mot f�rdragets bokstav och jag hoppas att det inte kommer till st�nd .
